module sequential_multiplier_rnl (clk,
    done,
    rst,
    start,
    multiplicand,
    multiplier,
    product);
 input clk;
 output done;
 input rst;
 input start;
 input [31:0] multiplicand;
 input [31:0] multiplier;
 output [63:0] product;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire \a[0] ;
 wire \a[10] ;
 wire \a[11] ;
 wire \a[12] ;
 wire \a[13] ;
 wire \a[14] ;
 wire \a[15] ;
 wire \a[16] ;
 wire \a[17] ;
 wire \a[18] ;
 wire \a[19] ;
 wire \a[1] ;
 wire \a[20] ;
 wire \a[21] ;
 wire \a[22] ;
 wire \a[23] ;
 wire \a[24] ;
 wire \a[25] ;
 wire \a[26] ;
 wire \a[27] ;
 wire \a[28] ;
 wire \a[29] ;
 wire \a[2] ;
 wire \a[30] ;
 wire \a[31] ;
 wire \a[3] ;
 wire \a[4] ;
 wire \a[5] ;
 wire \a[6] ;
 wire \a[7] ;
 wire \a[8] ;
 wire \a[9] ;
 wire \b[0] ;
 wire \b[10] ;
 wire \b[11] ;
 wire \b[12] ;
 wire \b[13] ;
 wire \b[14] ;
 wire \b[15] ;
 wire \b[16] ;
 wire \b[17] ;
 wire \b[18] ;
 wire \b[19] ;
 wire \b[1] ;
 wire \b[20] ;
 wire \b[21] ;
 wire \b[22] ;
 wire \b[23] ;
 wire \b[24] ;
 wire \b[25] ;
 wire \b[26] ;
 wire \b[27] ;
 wire \b[28] ;
 wire \b[29] ;
 wire \b[2] ;
 wire \b[30] ;
 wire \b[31] ;
 wire \b[3] ;
 wire \b[4] ;
 wire \b[5] ;
 wire \b[6] ;
 wire \b[7] ;
 wire \b[8] ;
 wire \b[9] ;
 wire \count[0] ;
 wire \count[1] ;
 wire \count[2] ;
 wire \count[3] ;
 wire \count[4] ;
 wire \count[5] ;
 wire \temp_product[0] ;
 wire \temp_product[10] ;
 wire \temp_product[11] ;
 wire \temp_product[12] ;
 wire \temp_product[13] ;
 wire \temp_product[14] ;
 wire \temp_product[15] ;
 wire \temp_product[16] ;
 wire \temp_product[17] ;
 wire \temp_product[18] ;
 wire \temp_product[19] ;
 wire \temp_product[1] ;
 wire \temp_product[20] ;
 wire \temp_product[21] ;
 wire \temp_product[22] ;
 wire \temp_product[23] ;
 wire \temp_product[24] ;
 wire \temp_product[25] ;
 wire \temp_product[26] ;
 wire \temp_product[27] ;
 wire \temp_product[28] ;
 wire \temp_product[29] ;
 wire \temp_product[2] ;
 wire \temp_product[30] ;
 wire \temp_product[31] ;
 wire \temp_product[32] ;
 wire \temp_product[33] ;
 wire \temp_product[34] ;
 wire \temp_product[35] ;
 wire \temp_product[36] ;
 wire \temp_product[37] ;
 wire \temp_product[38] ;
 wire \temp_product[39] ;
 wire \temp_product[3] ;
 wire \temp_product[40] ;
 wire \temp_product[41] ;
 wire \temp_product[42] ;
 wire \temp_product[43] ;
 wire \temp_product[44] ;
 wire \temp_product[45] ;
 wire \temp_product[46] ;
 wire \temp_product[47] ;
 wire \temp_product[48] ;
 wire \temp_product[49] ;
 wire \temp_product[4] ;
 wire \temp_product[50] ;
 wire \temp_product[51] ;
 wire \temp_product[52] ;
 wire \temp_product[53] ;
 wire \temp_product[54] ;
 wire \temp_product[55] ;
 wire \temp_product[56] ;
 wire \temp_product[57] ;
 wire \temp_product[58] ;
 wire \temp_product[59] ;
 wire \temp_product[5] ;
 wire \temp_product[60] ;
 wire \temp_product[61] ;
 wire \temp_product[62] ;
 wire \temp_product[63] ;
 wire \temp_product[6] ;
 wire \temp_product[7] ;
 wire \temp_product[8] ;
 wire \temp_product[9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;

 sky130_fd_sc_hd__inv_2 _0918_ (.A(net225),
    .Y(_0000_));
 sky130_fd_sc_hd__or2_1 _0919_ (.A(\count[1] ),
    .B(\count[0] ),
    .X(_0665_));
 sky130_fd_sc_hd__or2_1 _0920_ (.A(\count[2] ),
    .B(_0665_),
    .X(_0666_));
 sky130_fd_sc_hd__or2_1 _0921_ (.A(\count[3] ),
    .B(_0666_),
    .X(_0667_));
 sky130_fd_sc_hd__or2_1 _0922_ (.A(\count[4] ),
    .B(_0667_),
    .X(_0668_));
 sky130_fd_sc_hd__nor2_1 _0923_ (.A(\count[5] ),
    .B(_0668_),
    .Y(_0669_));
 sky130_fd_sc_hd__or2_1 _0924_ (.A(\count[5] ),
    .B(_0668_),
    .X(_0670_));
 sky130_fd_sc_hd__nor2_1 _0925_ (.A(net205),
    .B(_0670_),
    .Y(_0671_));
 sky130_fd_sc_hd__or2_1 _0926_ (.A(net203),
    .B(net182),
    .X(_0672_));
 sky130_fd_sc_hd__nor2_1 _0927_ (.A(net205),
    .B(net183),
    .Y(_0673_));
 sky130_fd_sc_hd__or2_2 _0928_ (.A(net203),
    .B(net183),
    .X(_0674_));
 sky130_fd_sc_hd__nor2_2 _0929_ (.A(\b[0] ),
    .B(_0674_),
    .Y(_0675_));
 sky130_fd_sc_hd__or2_1 _0930_ (.A(net181),
    .B(net152),
    .X(_0676_));
 sky130_fd_sc_hd__nand2_1 _0931_ (.A(\temp_product[31] ),
    .B(net191),
    .Y(_0677_));
 sky130_fd_sc_hd__or2_1 _0932_ (.A(\temp_product[31] ),
    .B(net191),
    .X(_0678_));
 sky130_fd_sc_hd__nand2_1 _0933_ (.A(_0677_),
    .B(_0678_),
    .Y(_0679_));
 sky130_fd_sc_hd__nand2_1 _0934_ (.A(\temp_product[30] ),
    .B(\a[30] ),
    .Y(_0680_));
 sky130_fd_sc_hd__or2_1 _0935_ (.A(\temp_product[30] ),
    .B(\a[30] ),
    .X(_0681_));
 sky130_fd_sc_hd__nand2_1 _0936_ (.A(_0680_),
    .B(_0681_),
    .Y(_0682_));
 sky130_fd_sc_hd__nor2_1 _0937_ (.A(\temp_product[29] ),
    .B(\a[29] ),
    .Y(_0683_));
 sky130_fd_sc_hd__and2_1 _0938_ (.A(\temp_product[29] ),
    .B(\a[29] ),
    .X(_0684_));
 sky130_fd_sc_hd__nand2_1 _0939_ (.A(\temp_product[28] ),
    .B(\a[28] ),
    .Y(_0685_));
 sky130_fd_sc_hd__and2b_1 _0940_ (.A_N(_0684_),
    .B(_0685_),
    .X(_0686_));
 sky130_fd_sc_hd__or2_1 _0941_ (.A(\temp_product[28] ),
    .B(\a[28] ),
    .X(_0687_));
 sky130_fd_sc_hd__nand2_1 _0942_ (.A(_0685_),
    .B(_0687_),
    .Y(_0688_));
 sky130_fd_sc_hd__nand2_1 _0943_ (.A(\temp_product[27] ),
    .B(\a[27] ),
    .Y(_0689_));
 sky130_fd_sc_hd__inv_2 _0944_ (.A(_0689_),
    .Y(_0690_));
 sky130_fd_sc_hd__nor2_1 _0945_ (.A(\temp_product[27] ),
    .B(\a[27] ),
    .Y(_0691_));
 sky130_fd_sc_hd__nand2_1 _0946_ (.A(\temp_product[26] ),
    .B(\a[26] ),
    .Y(_0692_));
 sky130_fd_sc_hd__a21o_1 _0947_ (.A1(_0689_),
    .A2(_0692_),
    .B1(_0691_),
    .X(_0693_));
 sky130_fd_sc_hd__or2_1 _0948_ (.A(_0690_),
    .B(_0691_),
    .X(_0694_));
 sky130_fd_sc_hd__or2_1 _0949_ (.A(\temp_product[26] ),
    .B(\a[26] ),
    .X(_0695_));
 sky130_fd_sc_hd__nand2_1 _0950_ (.A(_0692_),
    .B(_0695_),
    .Y(_0696_));
 sky130_fd_sc_hd__and2_1 _0951_ (.A(\temp_product[24] ),
    .B(\a[24] ),
    .X(_0697_));
 sky130_fd_sc_hd__a21o_1 _0952_ (.A1(\temp_product[25] ),
    .A2(\a[25] ),
    .B1(_0697_),
    .X(_0698_));
 sky130_fd_sc_hd__nor2_1 _0953_ (.A(\temp_product[24] ),
    .B(\a[24] ),
    .Y(_0699_));
 sky130_fd_sc_hd__nor2_1 _0954_ (.A(_0697_),
    .B(_0699_),
    .Y(_0700_));
 sky130_fd_sc_hd__and2_1 _0955_ (.A(\temp_product[23] ),
    .B(\a[23] ),
    .X(_0701_));
 sky130_fd_sc_hd__nand2_1 _0956_ (.A(\temp_product[22] ),
    .B(\a[22] ),
    .Y(_0702_));
 sky130_fd_sc_hd__nand2_1 _0957_ (.A(\temp_product[20] ),
    .B(\a[20] ),
    .Y(_0703_));
 sky130_fd_sc_hd__a22o_1 _0958_ (.A1(\temp_product[21] ),
    .A2(\a[21] ),
    .B1(\a[20] ),
    .B2(\temp_product[20] ),
    .X(_0704_));
 sky130_fd_sc_hd__inv_2 _0959_ (.A(_0704_),
    .Y(_0705_));
 sky130_fd_sc_hd__and2_1 _0960_ (.A(\temp_product[19] ),
    .B(\a[19] ),
    .X(_0706_));
 sky130_fd_sc_hd__nor2_1 _0961_ (.A(\temp_product[19] ),
    .B(\a[19] ),
    .Y(_0707_));
 sky130_fd_sc_hd__or2_1 _0962_ (.A(_0706_),
    .B(_0707_),
    .X(_0708_));
 sky130_fd_sc_hd__nand2_1 _0963_ (.A(\temp_product[18] ),
    .B(\a[18] ),
    .Y(_0709_));
 sky130_fd_sc_hd__or2_1 _0964_ (.A(\temp_product[18] ),
    .B(\a[18] ),
    .X(_0710_));
 sky130_fd_sc_hd__nand2_1 _0965_ (.A(_0709_),
    .B(_0710_),
    .Y(_0711_));
 sky130_fd_sc_hd__or2_1 _0966_ (.A(_0708_),
    .B(_0711_),
    .X(_0712_));
 sky130_fd_sc_hd__and2_1 _0967_ (.A(\temp_product[17] ),
    .B(\a[17] ),
    .X(_0713_));
 sky130_fd_sc_hd__nor2_1 _0968_ (.A(\temp_product[17] ),
    .B(\a[17] ),
    .Y(_0714_));
 sky130_fd_sc_hd__a21oi_1 _0969_ (.A1(\temp_product[16] ),
    .A2(\a[16] ),
    .B1(_0713_),
    .Y(_0715_));
 sky130_fd_sc_hd__nand2b_1 _0970_ (.A_N(_0706_),
    .B(_0709_),
    .Y(_0716_));
 sky130_fd_sc_hd__inv_2 _0971_ (.A(_0716_),
    .Y(_0717_));
 sky130_fd_sc_hd__o32a_1 _0972_ (.A1(_0712_),
    .A2(_0714_),
    .A3(_0715_),
    .B1(_0717_),
    .B2(_0707_),
    .X(_0718_));
 sky130_fd_sc_hd__or2_1 _0973_ (.A(\temp_product[20] ),
    .B(\a[20] ),
    .X(_0719_));
 sky130_fd_sc_hd__nor2_1 _0974_ (.A(\temp_product[23] ),
    .B(\a[23] ),
    .Y(_0720_));
 sky130_fd_sc_hd__or2_1 _0975_ (.A(\temp_product[22] ),
    .B(\a[22] ),
    .X(_0721_));
 sky130_fd_sc_hd__nand2_1 _0976_ (.A(_0703_),
    .B(_0719_),
    .Y(_0722_));
 sky130_fd_sc_hd__xnor2_1 _0977_ (.A(\temp_product[21] ),
    .B(\a[21] ),
    .Y(_0723_));
 sky130_fd_sc_hd__or2_1 _0978_ (.A(_0701_),
    .B(_0720_),
    .X(_0724_));
 sky130_fd_sc_hd__nand2_1 _0979_ (.A(_0702_),
    .B(_0721_),
    .Y(_0725_));
 sky130_fd_sc_hd__nor2_1 _0980_ (.A(_0724_),
    .B(_0725_),
    .Y(_0726_));
 sky130_fd_sc_hd__or4_1 _0981_ (.A(_0722_),
    .B(_0723_),
    .C(_0724_),
    .D(_0725_),
    .X(_0727_));
 sky130_fd_sc_hd__o22a_1 _0982_ (.A1(_0702_),
    .A2(_0720_),
    .B1(_0727_),
    .B2(_0718_),
    .X(_0728_));
 sky130_fd_sc_hd__o211a_1 _0983_ (.A1(\temp_product[21] ),
    .A2(\a[21] ),
    .B1(_0704_),
    .C1(_0726_),
    .X(_0729_));
 sky130_fd_sc_hd__or3b_1 _0984_ (.A(_0701_),
    .B(_0729_),
    .C_N(_0728_),
    .X(_0730_));
 sky130_fd_sc_hd__xnor2_1 _0985_ (.A(\temp_product[12] ),
    .B(\a[12] ),
    .Y(_0731_));
 sky130_fd_sc_hd__xnor2_1 _0986_ (.A(\temp_product[13] ),
    .B(\a[13] ),
    .Y(_0732_));
 sky130_fd_sc_hd__nand2_1 _0987_ (.A(\temp_product[14] ),
    .B(\a[14] ),
    .Y(_0733_));
 sky130_fd_sc_hd__or2_1 _0988_ (.A(\temp_product[14] ),
    .B(\a[14] ),
    .X(_0734_));
 sky130_fd_sc_hd__nand2_1 _0989_ (.A(_0733_),
    .B(_0734_),
    .Y(_0735_));
 sky130_fd_sc_hd__nand2_1 _0990_ (.A(\temp_product[15] ),
    .B(\a[15] ),
    .Y(_0736_));
 sky130_fd_sc_hd__or2_1 _0991_ (.A(\temp_product[15] ),
    .B(\a[15] ),
    .X(_0737_));
 sky130_fd_sc_hd__nand2_1 _0992_ (.A(_0736_),
    .B(_0737_),
    .Y(_0738_));
 sky130_fd_sc_hd__nor2_1 _0993_ (.A(_0735_),
    .B(_0738_),
    .Y(_0739_));
 sky130_fd_sc_hd__or4_1 _0994_ (.A(_0731_),
    .B(_0732_),
    .C(_0735_),
    .D(_0738_),
    .X(_0740_));
 sky130_fd_sc_hd__and2_1 _0995_ (.A(\temp_product[9] ),
    .B(\a[9] ),
    .X(_0741_));
 sky130_fd_sc_hd__nand2_1 _0996_ (.A(\temp_product[9] ),
    .B(\a[9] ),
    .Y(_0742_));
 sky130_fd_sc_hd__nand2_1 _0997_ (.A(\temp_product[8] ),
    .B(\a[8] ),
    .Y(_0743_));
 sky130_fd_sc_hd__nand2_1 _0998_ (.A(_0742_),
    .B(_0743_),
    .Y(_0744_));
 sky130_fd_sc_hd__xnor2_1 _0999_ (.A(\temp_product[11] ),
    .B(\a[11] ),
    .Y(_0745_));
 sky130_fd_sc_hd__nand2_1 _1000_ (.A(\temp_product[10] ),
    .B(\a[10] ),
    .Y(_0746_));
 sky130_fd_sc_hd__or2_1 _1001_ (.A(\temp_product[10] ),
    .B(\a[10] ),
    .X(_0747_));
 sky130_fd_sc_hd__nand2_1 _1002_ (.A(_0746_),
    .B(_0747_),
    .Y(_0748_));
 sky130_fd_sc_hd__nor2_1 _1003_ (.A(\temp_product[9] ),
    .B(\a[9] ),
    .Y(_0749_));
 sky130_fd_sc_hd__nor3_1 _1004_ (.A(_0745_),
    .B(_0748_),
    .C(_0749_),
    .Y(_0750_));
 sky130_fd_sc_hd__o211a_1 _1005_ (.A1(\temp_product[11] ),
    .A2(\a[11] ),
    .B1(\a[10] ),
    .C1(\temp_product[10] ),
    .X(_0751_));
 sky130_fd_sc_hd__a221o_1 _1006_ (.A1(\temp_product[11] ),
    .A2(\a[11] ),
    .B1(_0744_),
    .B2(_0750_),
    .C1(_0751_),
    .X(_0752_));
 sky130_fd_sc_hd__nor2_1 _1007_ (.A(\temp_product[3] ),
    .B(\a[3] ),
    .Y(_0753_));
 sky130_fd_sc_hd__nand2_1 _1008_ (.A(\temp_product[2] ),
    .B(\a[2] ),
    .Y(_0754_));
 sky130_fd_sc_hd__or2_1 _1009_ (.A(\temp_product[2] ),
    .B(\a[2] ),
    .X(_0755_));
 sky130_fd_sc_hd__nand2_1 _1010_ (.A(_0754_),
    .B(_0755_),
    .Y(_0756_));
 sky130_fd_sc_hd__nand2_1 _1011_ (.A(\temp_product[1] ),
    .B(\a[1] ),
    .Y(_0757_));
 sky130_fd_sc_hd__or2_1 _1012_ (.A(\temp_product[1] ),
    .B(\a[1] ),
    .X(_0758_));
 sky130_fd_sc_hd__nand4_1 _1013_ (.A(\temp_product[0] ),
    .B(\a[0] ),
    .C(_0757_),
    .D(_0758_),
    .Y(_0759_));
 sky130_fd_sc_hd__a21o_1 _1014_ (.A1(_0757_),
    .A2(_0759_),
    .B1(_0756_),
    .X(_0760_));
 sky130_fd_sc_hd__and2_1 _1015_ (.A(\temp_product[3] ),
    .B(\a[3] ),
    .X(_0761_));
 sky130_fd_sc_hd__nand2_1 _1016_ (.A(\temp_product[3] ),
    .B(\a[3] ),
    .Y(_0762_));
 sky130_fd_sc_hd__a31o_1 _1017_ (.A1(_0754_),
    .A2(_0760_),
    .A3(_0762_),
    .B1(_0753_),
    .X(_0763_));
 sky130_fd_sc_hd__or2_1 _1018_ (.A(\temp_product[7] ),
    .B(\a[7] ),
    .X(_0764_));
 sky130_fd_sc_hd__nand2_1 _1019_ (.A(\temp_product[7] ),
    .B(\a[7] ),
    .Y(_0765_));
 sky130_fd_sc_hd__xor2_1 _1020_ (.A(\temp_product[6] ),
    .B(\a[6] ),
    .X(_0766_));
 sky130_fd_sc_hd__nand3_1 _1021_ (.A(_0764_),
    .B(_0765_),
    .C(_0766_),
    .Y(_0767_));
 sky130_fd_sc_hd__xnor2_1 _1022_ (.A(\temp_product[4] ),
    .B(\a[4] ),
    .Y(_0768_));
 sky130_fd_sc_hd__and2_1 _1023_ (.A(\temp_product[5] ),
    .B(\a[5] ),
    .X(_0769_));
 sky130_fd_sc_hd__nor2_1 _1024_ (.A(\temp_product[5] ),
    .B(\a[5] ),
    .Y(_0770_));
 sky130_fd_sc_hd__nor2_1 _1025_ (.A(_0769_),
    .B(_0770_),
    .Y(_0771_));
 sky130_fd_sc_hd__or3b_1 _1026_ (.A(_0767_),
    .B(_0768_),
    .C_N(_0771_),
    .X(_0772_));
 sky130_fd_sc_hd__a311o_1 _1027_ (.A1(_0754_),
    .A2(_0760_),
    .A3(_0762_),
    .B1(_0772_),
    .C1(_0753_),
    .X(_0773_));
 sky130_fd_sc_hd__a21o_1 _1028_ (.A1(\temp_product[4] ),
    .A2(\a[4] ),
    .B1(_0769_),
    .X(_0774_));
 sky130_fd_sc_hd__nand2b_1 _1029_ (.A_N(_0770_),
    .B(_0774_),
    .Y(_0775_));
 sky130_fd_sc_hd__a22o_1 _1030_ (.A1(\temp_product[7] ),
    .A2(\a[7] ),
    .B1(\a[6] ),
    .B2(\temp_product[6] ),
    .X(_0776_));
 sky130_fd_sc_hd__o2bb2a_1 _1031_ (.A1_N(_0764_),
    .A2_N(_0776_),
    .B1(_0775_),
    .B2(_0767_),
    .X(_0777_));
 sky130_fd_sc_hd__or2_1 _1032_ (.A(\temp_product[8] ),
    .B(\a[8] ),
    .X(_0778_));
 sky130_fd_sc_hd__nand2_1 _1033_ (.A(_0743_),
    .B(_0778_),
    .Y(_0779_));
 sky130_fd_sc_hd__nand2_1 _1034_ (.A(_0742_),
    .B(_0750_),
    .Y(_0780_));
 sky130_fd_sc_hd__a21o_1 _1035_ (.A1(_0773_),
    .A2(_0777_),
    .B1(_0779_),
    .X(_0781_));
 sky130_fd_sc_hd__o21ba_1 _1036_ (.A1(_0780_),
    .A2(_0781_),
    .B1_N(_0752_),
    .X(_0782_));
 sky130_fd_sc_hd__a22o_1 _1037_ (.A1(\temp_product[13] ),
    .A2(\a[13] ),
    .B1(\a[12] ),
    .B2(\temp_product[12] ),
    .X(_0783_));
 sky130_fd_sc_hd__o211a_1 _1038_ (.A1(\temp_product[13] ),
    .A2(\a[13] ),
    .B1(_0739_),
    .C1(_0783_),
    .X(_0784_));
 sky130_fd_sc_hd__a31oi_2 _1039_ (.A1(\temp_product[14] ),
    .A2(\a[14] ),
    .A3(_0737_),
    .B1(_0784_),
    .Y(_0785_));
 sky130_fd_sc_hd__o211ai_4 _1040_ (.A1(_0740_),
    .A2(_0782_),
    .B1(_0785_),
    .C1(_0736_),
    .Y(_0786_));
 sky130_fd_sc_hd__xor2_1 _1041_ (.A(\temp_product[16] ),
    .B(\a[16] ),
    .X(_0787_));
 sky130_fd_sc_hd__nor2_1 _1042_ (.A(_0713_),
    .B(_0714_),
    .Y(_0788_));
 sky130_fd_sc_hd__and4bb_1 _1043_ (.A_N(_0712_),
    .B_N(_0727_),
    .C(_0787_),
    .D(_0788_),
    .X(_0789_));
 sky130_fd_sc_hd__and2_1 _1044_ (.A(_0786_),
    .B(_0789_),
    .X(_0790_));
 sky130_fd_sc_hd__o21a_1 _1045_ (.A1(_0730_),
    .A2(_0790_),
    .B1(_0700_),
    .X(_0791_));
 sky130_fd_sc_hd__o22a_1 _1046_ (.A1(\temp_product[25] ),
    .A2(\a[25] ),
    .B1(_0698_),
    .B2(_0791_),
    .X(_0792_));
 sky130_fd_sc_hd__or3b_1 _1047_ (.A(_0694_),
    .B(_0696_),
    .C_N(_0792_),
    .X(_0793_));
 sky130_fd_sc_hd__a21o_1 _1048_ (.A1(_0693_),
    .A2(_0793_),
    .B1(_0688_),
    .X(_0794_));
 sky130_fd_sc_hd__a21o_1 _1049_ (.A1(_0686_),
    .A2(_0794_),
    .B1(_0683_),
    .X(_0795_));
 sky130_fd_sc_hd__or2_1 _1050_ (.A(_0682_),
    .B(_0795_),
    .X(_0796_));
 sky130_fd_sc_hd__nand3_1 _1051_ (.A(_0679_),
    .B(_0680_),
    .C(_0796_),
    .Y(_0797_));
 sky130_fd_sc_hd__and2_1 _1052_ (.A(\b[0] ),
    .B(net159),
    .X(_0798_));
 sky130_fd_sc_hd__a21o_1 _1053_ (.A1(_0680_),
    .A2(_0796_),
    .B1(_0679_),
    .X(_0799_));
 sky130_fd_sc_hd__a32o_1 _1054_ (.A1(_0797_),
    .A2(net144),
    .A3(_0799_),
    .B1(net133),
    .B2(\temp_product[31] ),
    .X(_0397_));
 sky130_fd_sc_hd__nand2_1 _1055_ (.A(_0682_),
    .B(_0795_),
    .Y(_0800_));
 sky130_fd_sc_hd__a32o_1 _1056_ (.A1(_0796_),
    .A2(net147),
    .A3(_0800_),
    .B1(net133),
    .B2(\temp_product[30] ),
    .X(_0396_));
 sky130_fd_sc_hd__or2_1 _1057_ (.A(_0683_),
    .B(_0684_),
    .X(_0801_));
 sky130_fd_sc_hd__a21o_1 _1058_ (.A1(_0685_),
    .A2(_0794_),
    .B1(_0801_),
    .X(_0802_));
 sky130_fd_sc_hd__nand3_1 _1059_ (.A(_0685_),
    .B(_0794_),
    .C(_0801_),
    .Y(_0803_));
 sky130_fd_sc_hd__a32o_1 _1060_ (.A1(net147),
    .A2(_0802_),
    .A3(_0803_),
    .B1(net133),
    .B2(\temp_product[29] ),
    .X(_0395_));
 sky130_fd_sc_hd__nand3_1 _1061_ (.A(_0688_),
    .B(_0693_),
    .C(_0793_),
    .Y(_0804_));
 sky130_fd_sc_hd__a32o_1 _1062_ (.A1(_0794_),
    .A2(net147),
    .A3(_0804_),
    .B1(net133),
    .B2(\temp_product[28] ),
    .X(_0394_));
 sky130_fd_sc_hd__a21bo_1 _1063_ (.A1(_0695_),
    .A2(_0792_),
    .B1_N(_0692_),
    .X(_0805_));
 sky130_fd_sc_hd__xnor2_1 _1064_ (.A(_0694_),
    .B(_0805_),
    .Y(_0806_));
 sky130_fd_sc_hd__a22o_1 _1065_ (.A1(\temp_product[27] ),
    .A2(net132),
    .B1(net144),
    .B2(_0806_),
    .X(_0393_));
 sky130_fd_sc_hd__xnor2_1 _1066_ (.A(_0696_),
    .B(_0792_),
    .Y(_0807_));
 sky130_fd_sc_hd__a22o_1 _1067_ (.A1(\temp_product[26] ),
    .A2(net135),
    .B1(net146),
    .B2(_0807_),
    .X(_0392_));
 sky130_fd_sc_hd__xor2_1 _1068_ (.A(\temp_product[25] ),
    .B(\a[25] ),
    .X(_0808_));
 sky130_fd_sc_hd__o21ai_1 _1069_ (.A1(_0697_),
    .A2(_0791_),
    .B1(_0808_),
    .Y(_0809_));
 sky130_fd_sc_hd__or3_1 _1070_ (.A(_0697_),
    .B(_0791_),
    .C(_0808_),
    .X(_0810_));
 sky130_fd_sc_hd__a32o_1 _1071_ (.A1(net146),
    .A2(_0809_),
    .A3(_0810_),
    .B1(net135),
    .B2(\temp_product[25] ),
    .X(_0391_));
 sky130_fd_sc_hd__or3_1 _1072_ (.A(_0700_),
    .B(_0730_),
    .C(_0790_),
    .X(_0811_));
 sky130_fd_sc_hd__and2b_1 _1073_ (.A_N(_0791_),
    .B(net146),
    .X(_0812_));
 sky130_fd_sc_hd__a22o_1 _1074_ (.A1(\temp_product[24] ),
    .A2(net135),
    .B1(_0811_),
    .B2(_0812_),
    .X(_0390_));
 sky130_fd_sc_hd__nand2_1 _1075_ (.A(_0786_),
    .B(_0787_),
    .Y(_0813_));
 sky130_fd_sc_hd__a22o_1 _1076_ (.A1(\temp_product[16] ),
    .A2(\a[16] ),
    .B1(_0786_),
    .B2(_0787_),
    .X(_0814_));
 sky130_fd_sc_hd__o21bai_1 _1077_ (.A1(_0713_),
    .A2(_0814_),
    .B1_N(_0714_),
    .Y(_0815_));
 sky130_fd_sc_hd__or2_1 _1078_ (.A(_0711_),
    .B(_0815_),
    .X(_0816_));
 sky130_fd_sc_hd__a211o_1 _1079_ (.A1(_0717_),
    .A2(_0816_),
    .B1(_0722_),
    .C1(_0707_),
    .X(_0817_));
 sky130_fd_sc_hd__a2bb2o_1 _1080_ (.A1_N(\temp_product[21] ),
    .A2_N(\a[21] ),
    .B1(_0705_),
    .B2(_0817_),
    .X(_0818_));
 sky130_fd_sc_hd__or2_1 _1081_ (.A(_0725_),
    .B(_0818_),
    .X(_0819_));
 sky130_fd_sc_hd__nand3_1 _1082_ (.A(_0702_),
    .B(_0724_),
    .C(_0819_),
    .Y(_0820_));
 sky130_fd_sc_hd__a21o_1 _1083_ (.A1(_0702_),
    .A2(_0819_),
    .B1(_0724_),
    .X(_0821_));
 sky130_fd_sc_hd__a32o_1 _1084_ (.A1(net146),
    .A2(_0820_),
    .A3(_0821_),
    .B1(net135),
    .B2(\temp_product[23] ),
    .X(_0389_));
 sky130_fd_sc_hd__nand2_1 _1085_ (.A(_0725_),
    .B(_0818_),
    .Y(_0822_));
 sky130_fd_sc_hd__a32o_1 _1086_ (.A1(net146),
    .A2(_0819_),
    .A3(_0822_),
    .B1(net135),
    .B2(\temp_product[22] ),
    .X(_0388_));
 sky130_fd_sc_hd__nand3_1 _1087_ (.A(_0703_),
    .B(_0723_),
    .C(_0817_),
    .Y(_0823_));
 sky130_fd_sc_hd__a21o_1 _1088_ (.A1(_0703_),
    .A2(_0817_),
    .B1(_0723_),
    .X(_0824_));
 sky130_fd_sc_hd__a32o_1 _1089_ (.A1(net146),
    .A2(_0823_),
    .A3(_0824_),
    .B1(net135),
    .B2(\temp_product[21] ),
    .X(_0387_));
 sky130_fd_sc_hd__o221ai_1 _1090_ (.A1(_0707_),
    .A2(_0717_),
    .B1(_0815_),
    .B2(_0712_),
    .C1(_0722_),
    .Y(_0825_));
 sky130_fd_sc_hd__a32o_1 _1091_ (.A1(net146),
    .A2(_0817_),
    .A3(_0825_),
    .B1(net135),
    .B2(\temp_product[20] ),
    .X(_0386_));
 sky130_fd_sc_hd__nand2_1 _1092_ (.A(_0709_),
    .B(_0816_),
    .Y(_0826_));
 sky130_fd_sc_hd__xnor2_1 _1093_ (.A(_0708_),
    .B(_0826_),
    .Y(_0827_));
 sky130_fd_sc_hd__a22o_1 _1094_ (.A1(\temp_product[19] ),
    .A2(net134),
    .B1(net145),
    .B2(_0827_),
    .X(_0385_));
 sky130_fd_sc_hd__nand2_1 _1095_ (.A(_0711_),
    .B(_0815_),
    .Y(_0828_));
 sky130_fd_sc_hd__a32o_1 _1096_ (.A1(net145),
    .A2(_0816_),
    .A3(_0828_),
    .B1(net134),
    .B2(\temp_product[18] ),
    .X(_0384_));
 sky130_fd_sc_hd__xor2_1 _1097_ (.A(_0788_),
    .B(_0814_),
    .X(_0829_));
 sky130_fd_sc_hd__a22o_1 _1098_ (.A1(\temp_product[17] ),
    .A2(net134),
    .B1(net145),
    .B2(_0829_),
    .X(_0383_));
 sky130_fd_sc_hd__or2_1 _1099_ (.A(_0786_),
    .B(_0787_),
    .X(_0830_));
 sky130_fd_sc_hd__a32o_1 _1100_ (.A1(net145),
    .A2(_0813_),
    .A3(_0830_),
    .B1(net134),
    .B2(\temp_product[16] ),
    .X(_0382_));
 sky130_fd_sc_hd__nor2_1 _1101_ (.A(_0731_),
    .B(_0782_),
    .Y(_0831_));
 sky130_fd_sc_hd__or2_1 _1102_ (.A(_0731_),
    .B(_0782_),
    .X(_0832_));
 sky130_fd_sc_hd__o22a_1 _1103_ (.A1(\temp_product[13] ),
    .A2(\a[13] ),
    .B1(_0783_),
    .B2(_0831_),
    .X(_0833_));
 sky130_fd_sc_hd__a21bo_1 _1104_ (.A1(_0734_),
    .A2(_0833_),
    .B1_N(_0733_),
    .X(_0834_));
 sky130_fd_sc_hd__xnor2_1 _1105_ (.A(_0738_),
    .B(_0834_),
    .Y(_0835_));
 sky130_fd_sc_hd__a22o_1 _1106_ (.A1(\temp_product[15] ),
    .A2(net134),
    .B1(net145),
    .B2(_0835_),
    .X(_0381_));
 sky130_fd_sc_hd__xnor2_1 _1107_ (.A(_0735_),
    .B(_0833_),
    .Y(_0836_));
 sky130_fd_sc_hd__a22o_1 _1108_ (.A1(\temp_product[14] ),
    .A2(net134),
    .B1(net145),
    .B2(_0836_),
    .X(_0380_));
 sky130_fd_sc_hd__a21o_1 _1109_ (.A1(\temp_product[12] ),
    .A2(\a[12] ),
    .B1(_0831_),
    .X(_0837_));
 sky130_fd_sc_hd__xnor2_1 _1110_ (.A(_0732_),
    .B(_0837_),
    .Y(_0838_));
 sky130_fd_sc_hd__a22o_1 _1111_ (.A1(\temp_product[13] ),
    .A2(net134),
    .B1(net145),
    .B2(_0838_),
    .X(_0379_));
 sky130_fd_sc_hd__nand2_1 _1112_ (.A(_0731_),
    .B(_0782_),
    .Y(_0839_));
 sky130_fd_sc_hd__a32o_1 _1113_ (.A1(net145),
    .A2(_0832_),
    .A3(_0839_),
    .B1(net134),
    .B2(\temp_product[12] ),
    .X(_0378_));
 sky130_fd_sc_hd__a31o_1 _1114_ (.A1(_0742_),
    .A2(_0743_),
    .A3(_0781_),
    .B1(_0749_),
    .X(_0840_));
 sky130_fd_sc_hd__or2_1 _1115_ (.A(_0748_),
    .B(_0840_),
    .X(_0841_));
 sky130_fd_sc_hd__nand3_1 _1116_ (.A(_0745_),
    .B(_0746_),
    .C(_0841_),
    .Y(_0842_));
 sky130_fd_sc_hd__a21o_1 _1117_ (.A1(_0746_),
    .A2(_0841_),
    .B1(_0745_),
    .X(_0843_));
 sky130_fd_sc_hd__a32o_1 _1118_ (.A1(net145),
    .A2(_0842_),
    .A3(_0843_),
    .B1(net134),
    .B2(\temp_product[11] ),
    .X(_0377_));
 sky130_fd_sc_hd__nand2_1 _1119_ (.A(_0748_),
    .B(_0840_),
    .Y(_0844_));
 sky130_fd_sc_hd__a32o_1 _1120_ (.A1(net145),
    .A2(_0841_),
    .A3(_0844_),
    .B1(net134),
    .B2(\temp_product[10] ),
    .X(_0376_));
 sky130_fd_sc_hd__a211o_1 _1121_ (.A1(_0743_),
    .A2(_0781_),
    .B1(_0749_),
    .C1(_0741_),
    .X(_0845_));
 sky130_fd_sc_hd__o211ai_1 _1122_ (.A1(_0741_),
    .A2(_0749_),
    .B1(_0781_),
    .C1(_0743_),
    .Y(_0846_));
 sky130_fd_sc_hd__a32o_1 _1123_ (.A1(net144),
    .A2(_0845_),
    .A3(_0846_),
    .B1(net132),
    .B2(\temp_product[9] ),
    .X(_0375_));
 sky130_fd_sc_hd__and3_1 _1124_ (.A(_0773_),
    .B(_0777_),
    .C(_0779_),
    .X(_0847_));
 sky130_fd_sc_hd__nand2_1 _1125_ (.A(_0781_),
    .B(net144),
    .Y(_0848_));
 sky130_fd_sc_hd__a2bb2o_1 _1126_ (.A1_N(_0847_),
    .A2_N(_0848_),
    .B1(\temp_product[8] ),
    .B2(net132),
    .X(_0374_));
 sky130_fd_sc_hd__nor2_1 _1127_ (.A(_0763_),
    .B(_0768_),
    .Y(_0849_));
 sky130_fd_sc_hd__o21ba_1 _1128_ (.A1(_0774_),
    .A2(_0849_),
    .B1_N(_0770_),
    .X(_0850_));
 sky130_fd_sc_hd__and2_1 _1129_ (.A(_0766_),
    .B(_0850_),
    .X(_0851_));
 sky130_fd_sc_hd__a21o_1 _1130_ (.A1(\temp_product[6] ),
    .A2(\a[6] ),
    .B1(_0851_),
    .X(_0852_));
 sky130_fd_sc_hd__a21o_1 _1131_ (.A1(_0764_),
    .A2(_0765_),
    .B1(_0852_),
    .X(_0853_));
 sky130_fd_sc_hd__nand3_1 _1132_ (.A(_0764_),
    .B(_0765_),
    .C(_0852_),
    .Y(_0854_));
 sky130_fd_sc_hd__a32o_1 _1133_ (.A1(net144),
    .A2(_0853_),
    .A3(_0854_),
    .B1(net132),
    .B2(\temp_product[7] ),
    .X(_0373_));
 sky130_fd_sc_hd__nor2_1 _1134_ (.A(_0766_),
    .B(_0850_),
    .Y(_0855_));
 sky130_fd_sc_hd__nor2_1 _1135_ (.A(_0851_),
    .B(_0855_),
    .Y(_0856_));
 sky130_fd_sc_hd__a22o_1 _1136_ (.A1(\temp_product[6] ),
    .A2(net132),
    .B1(net144),
    .B2(_0856_),
    .X(_0372_));
 sky130_fd_sc_hd__a21oi_1 _1137_ (.A1(\temp_product[4] ),
    .A2(\a[4] ),
    .B1(_0849_),
    .Y(_0857_));
 sky130_fd_sc_hd__xnor2_1 _1138_ (.A(_0771_),
    .B(_0857_),
    .Y(_0858_));
 sky130_fd_sc_hd__a22o_1 _1139_ (.A1(\temp_product[5] ),
    .A2(net132),
    .B1(net144),
    .B2(_0858_),
    .X(_0371_));
 sky130_fd_sc_hd__nand2_1 _1140_ (.A(_0763_),
    .B(_0768_),
    .Y(_0859_));
 sky130_fd_sc_hd__and3b_1 _1141_ (.A_N(_0849_),
    .B(_0859_),
    .C(net144),
    .X(_0860_));
 sky130_fd_sc_hd__a21o_1 _1142_ (.A1(\temp_product[4] ),
    .A2(net132),
    .B1(_0860_),
    .X(_0370_));
 sky130_fd_sc_hd__a211o_1 _1143_ (.A1(_0754_),
    .A2(_0760_),
    .B1(_0761_),
    .C1(_0753_),
    .X(_0861_));
 sky130_fd_sc_hd__o211ai_1 _1144_ (.A1(_0753_),
    .A2(_0761_),
    .B1(_0760_),
    .C1(_0754_),
    .Y(_0862_));
 sky130_fd_sc_hd__a32o_1 _1145_ (.A1(net144),
    .A2(_0861_),
    .A3(_0862_),
    .B1(net132),
    .B2(\temp_product[3] ),
    .X(_0369_));
 sky130_fd_sc_hd__nand3_1 _1146_ (.A(_0756_),
    .B(_0757_),
    .C(_0759_),
    .Y(_0863_));
 sky130_fd_sc_hd__a32o_1 _1147_ (.A1(_0760_),
    .A2(net144),
    .A3(_0863_),
    .B1(net133),
    .B2(\temp_product[2] ),
    .X(_0368_));
 sky130_fd_sc_hd__a22o_1 _1148_ (.A1(\temp_product[0] ),
    .A2(\a[0] ),
    .B1(_0757_),
    .B2(_0758_),
    .X(_0864_));
 sky130_fd_sc_hd__a32o_1 _1149_ (.A1(_0759_),
    .A2(net147),
    .A3(_0864_),
    .B1(net132),
    .B2(\temp_product[1] ),
    .X(_0367_));
 sky130_fd_sc_hd__o211a_1 _1150_ (.A1(\b[0] ),
    .A2(_0674_),
    .B1(net168),
    .C1(\a[0] ),
    .X(_0865_));
 sky130_fd_sc_hd__a21oi_1 _1151_ (.A1(\temp_product[0] ),
    .A2(\a[0] ),
    .B1(net202),
    .Y(_0866_));
 sky130_fd_sc_hd__o22a_1 _1152_ (.A1(\temp_product[0] ),
    .A2(_0865_),
    .B1(_0866_),
    .B2(net132),
    .X(_0366_));
 sky130_fd_sc_hd__mux2_1 _1153_ (.A0(\b[31] ),
    .A1(net56),
    .S(net202),
    .X(_0867_));
 sky130_fd_sc_hd__mux2_1 _1154_ (.A0(\b[30] ),
    .A1(_0867_),
    .S(net168),
    .X(_0365_));
 sky130_fd_sc_hd__and2_1 _1155_ (.A(net202),
    .B(net54),
    .X(_0868_));
 sky130_fd_sc_hd__a221o_1 _1156_ (.A1(\b[29] ),
    .A2(net177),
    .B1(net160),
    .B2(\b[30] ),
    .C1(_0868_),
    .X(_0364_));
 sky130_fd_sc_hd__and2_1 _1157_ (.A(net202),
    .B(net53),
    .X(_0869_));
 sky130_fd_sc_hd__a221o_1 _1158_ (.A1(\b[28] ),
    .A2(net177),
    .B1(net160),
    .B2(\b[29] ),
    .C1(_0869_),
    .X(_0363_));
 sky130_fd_sc_hd__and2_1 _1159_ (.A(net203),
    .B(net52),
    .X(_0870_));
 sky130_fd_sc_hd__a221o_1 _1160_ (.A1(\b[27] ),
    .A2(net177),
    .B1(net160),
    .B2(\b[28] ),
    .C1(_0870_),
    .X(_0362_));
 sky130_fd_sc_hd__and2_1 _1161_ (.A(net203),
    .B(net51),
    .X(_0871_));
 sky130_fd_sc_hd__a221o_1 _1162_ (.A1(\b[26] ),
    .A2(net177),
    .B1(net160),
    .B2(\b[27] ),
    .C1(_0871_),
    .X(_0361_));
 sky130_fd_sc_hd__and2_1 _1163_ (.A(net203),
    .B(net50),
    .X(_0872_));
 sky130_fd_sc_hd__a221o_1 _1164_ (.A1(\b[25] ),
    .A2(net177),
    .B1(net160),
    .B2(\b[26] ),
    .C1(_0872_),
    .X(_0360_));
 sky130_fd_sc_hd__and2_1 _1165_ (.A(net204),
    .B(net49),
    .X(_0873_));
 sky130_fd_sc_hd__a221o_1 _1166_ (.A1(\b[24] ),
    .A2(net177),
    .B1(net160),
    .B2(\b[25] ),
    .C1(_0873_),
    .X(_0359_));
 sky130_fd_sc_hd__and2_1 _1167_ (.A(net204),
    .B(net48),
    .X(_0874_));
 sky130_fd_sc_hd__a221o_1 _1168_ (.A1(\b[23] ),
    .A2(net176),
    .B1(net159),
    .B2(\b[24] ),
    .C1(_0874_),
    .X(_0358_));
 sky130_fd_sc_hd__and2_1 _1169_ (.A(net202),
    .B(net47),
    .X(_0875_));
 sky130_fd_sc_hd__a221o_1 _1170_ (.A1(\b[22] ),
    .A2(net176),
    .B1(net159),
    .B2(\b[23] ),
    .C1(_0875_),
    .X(_0357_));
 sky130_fd_sc_hd__and2_1 _1171_ (.A(net202),
    .B(net46),
    .X(_0876_));
 sky130_fd_sc_hd__a221o_1 _1172_ (.A1(\b[21] ),
    .A2(net176),
    .B1(net159),
    .B2(\b[22] ),
    .C1(_0876_),
    .X(_0356_));
 sky130_fd_sc_hd__and2_1 _1173_ (.A(net202),
    .B(net45),
    .X(_0877_));
 sky130_fd_sc_hd__a221o_1 _1174_ (.A1(\b[20] ),
    .A2(net176),
    .B1(net159),
    .B2(\b[21] ),
    .C1(_0877_),
    .X(_0355_));
 sky130_fd_sc_hd__and2_1 _1175_ (.A(net199),
    .B(net43),
    .X(_0878_));
 sky130_fd_sc_hd__a221o_1 _1176_ (.A1(\b[19] ),
    .A2(net176),
    .B1(net159),
    .B2(\b[20] ),
    .C1(_0878_),
    .X(_0354_));
 sky130_fd_sc_hd__and2_1 _1177_ (.A(net199),
    .B(net42),
    .X(_0879_));
 sky130_fd_sc_hd__a221o_1 _1178_ (.A1(\b[18] ),
    .A2(net175),
    .B1(net158),
    .B2(\b[19] ),
    .C1(_0879_),
    .X(_0353_));
 sky130_fd_sc_hd__and2_1 _1179_ (.A(net199),
    .B(net41),
    .X(_0880_));
 sky130_fd_sc_hd__a221o_1 _1180_ (.A1(\b[17] ),
    .A2(net174),
    .B1(net157),
    .B2(\b[18] ),
    .C1(_0880_),
    .X(_0352_));
 sky130_fd_sc_hd__and2_1 _1181_ (.A(net199),
    .B(net40),
    .X(_0881_));
 sky130_fd_sc_hd__a221o_1 _1182_ (.A1(\b[16] ),
    .A2(net174),
    .B1(net157),
    .B2(\b[17] ),
    .C1(_0881_),
    .X(_0351_));
 sky130_fd_sc_hd__and2_1 _1183_ (.A(net197),
    .B(net39),
    .X(_0882_));
 sky130_fd_sc_hd__a221o_1 _1184_ (.A1(\b[15] ),
    .A2(net174),
    .B1(net157),
    .B2(\b[16] ),
    .C1(_0882_),
    .X(_0350_));
 sky130_fd_sc_hd__and2_1 _1185_ (.A(net196),
    .B(net38),
    .X(_0883_));
 sky130_fd_sc_hd__a221o_1 _1186_ (.A1(\b[14] ),
    .A2(net173),
    .B1(net156),
    .B2(\b[15] ),
    .C1(_0883_),
    .X(_0349_));
 sky130_fd_sc_hd__and2_1 _1187_ (.A(net196),
    .B(net37),
    .X(_0884_));
 sky130_fd_sc_hd__a221o_1 _1188_ (.A1(\b[13] ),
    .A2(net173),
    .B1(net156),
    .B2(\b[14] ),
    .C1(_0884_),
    .X(_0348_));
 sky130_fd_sc_hd__and2_1 _1189_ (.A(net196),
    .B(net36),
    .X(_0885_));
 sky130_fd_sc_hd__a221o_1 _1190_ (.A1(\b[12] ),
    .A2(net173),
    .B1(net156),
    .B2(\b[13] ),
    .C1(_0885_),
    .X(_0347_));
 sky130_fd_sc_hd__and2_1 _1191_ (.A(net196),
    .B(net35),
    .X(_0886_));
 sky130_fd_sc_hd__a221o_1 _1192_ (.A1(\b[11] ),
    .A2(net173),
    .B1(net156),
    .B2(\b[12] ),
    .C1(_0886_),
    .X(_0346_));
 sky130_fd_sc_hd__and2_1 _1193_ (.A(net197),
    .B(net34),
    .X(_0887_));
 sky130_fd_sc_hd__a221o_1 _1194_ (.A1(\b[10] ),
    .A2(net173),
    .B1(net156),
    .B2(\b[11] ),
    .C1(_0887_),
    .X(_0345_));
 sky130_fd_sc_hd__and2_1 _1195_ (.A(net197),
    .B(net64),
    .X(_0888_));
 sky130_fd_sc_hd__a221o_1 _1196_ (.A1(\b[9] ),
    .A2(net173),
    .B1(net156),
    .B2(\b[10] ),
    .C1(_0888_),
    .X(_0344_));
 sky130_fd_sc_hd__and2_1 _1197_ (.A(net197),
    .B(net63),
    .X(_0889_));
 sky130_fd_sc_hd__a221o_1 _1198_ (.A1(\b[8] ),
    .A2(net173),
    .B1(net156),
    .B2(\b[9] ),
    .C1(_0889_),
    .X(_0343_));
 sky130_fd_sc_hd__and2_1 _1199_ (.A(net199),
    .B(net62),
    .X(_0890_));
 sky130_fd_sc_hd__a221o_1 _1200_ (.A1(\b[7] ),
    .A2(net174),
    .B1(net157),
    .B2(\b[8] ),
    .C1(_0890_),
    .X(_0342_));
 sky130_fd_sc_hd__and2_1 _1201_ (.A(net199),
    .B(net61),
    .X(_0891_));
 sky130_fd_sc_hd__a221o_1 _1202_ (.A1(\b[6] ),
    .A2(net174),
    .B1(net157),
    .B2(\b[7] ),
    .C1(_0891_),
    .X(_0341_));
 sky130_fd_sc_hd__and2_1 _1203_ (.A(net197),
    .B(net60),
    .X(_0892_));
 sky130_fd_sc_hd__a221o_1 _1204_ (.A1(\b[5] ),
    .A2(net174),
    .B1(net157),
    .B2(\b[6] ),
    .C1(_0892_),
    .X(_0340_));
 sky130_fd_sc_hd__and2_1 _1205_ (.A(net199),
    .B(net59),
    .X(_0893_));
 sky130_fd_sc_hd__a221o_1 _1206_ (.A1(\b[4] ),
    .A2(net176),
    .B1(net159),
    .B2(\b[5] ),
    .C1(_0893_),
    .X(_0339_));
 sky130_fd_sc_hd__and2_1 _1207_ (.A(net204),
    .B(net58),
    .X(_0894_));
 sky130_fd_sc_hd__a221o_1 _1208_ (.A1(\b[3] ),
    .A2(net177),
    .B1(net160),
    .B2(\b[4] ),
    .C1(_0894_),
    .X(_0338_));
 sky130_fd_sc_hd__and2_1 _1209_ (.A(net204),
    .B(net55),
    .X(_0895_));
 sky130_fd_sc_hd__a221o_1 _1210_ (.A1(\b[2] ),
    .A2(net176),
    .B1(net159),
    .B2(\b[3] ),
    .C1(_0895_),
    .X(_0337_));
 sky130_fd_sc_hd__and2_1 _1211_ (.A(net204),
    .B(net44),
    .X(_0896_));
 sky130_fd_sc_hd__a221o_1 _1212_ (.A1(\b[1] ),
    .A2(net176),
    .B1(net159),
    .B2(\b[2] ),
    .C1(_0896_),
    .X(_0336_));
 sky130_fd_sc_hd__and2_1 _1213_ (.A(net202),
    .B(net33),
    .X(_0897_));
 sky130_fd_sc_hd__a221o_1 _1214_ (.A1(\b[0] ),
    .A2(net176),
    .B1(net159),
    .B2(\b[1] ),
    .C1(_0897_),
    .X(_0335_));
 sky130_fd_sc_hd__and2_1 _1215_ (.A(net203),
    .B(net25),
    .X(_0898_));
 sky130_fd_sc_hd__a221o_1 _1216_ (.A1(net191),
    .A2(net178),
    .B1(net161),
    .B2(\a[30] ),
    .C1(_0898_),
    .X(_0334_));
 sky130_fd_sc_hd__and2_1 _1217_ (.A(net204),
    .B(net24),
    .X(_0899_));
 sky130_fd_sc_hd__a221o_1 _1218_ (.A1(\a[30] ),
    .A2(net178),
    .B1(net161),
    .B2(\a[29] ),
    .C1(_0899_),
    .X(_0333_));
 sky130_fd_sc_hd__and2_1 _1219_ (.A(net196),
    .B(net22),
    .X(_0900_));
 sky130_fd_sc_hd__a221o_1 _1220_ (.A1(\a[29] ),
    .A2(net175),
    .B1(net158),
    .B2(\a[28] ),
    .C1(_0900_),
    .X(_0332_));
 sky130_fd_sc_hd__and2_1 _1221_ (.A(net199),
    .B(net21),
    .X(_0901_));
 sky130_fd_sc_hd__a221o_1 _1222_ (.A1(\a[28] ),
    .A2(net175),
    .B1(net158),
    .B2(\a[27] ),
    .C1(_0901_),
    .X(_0331_));
 sky130_fd_sc_hd__and2_1 _1223_ (.A(net198),
    .B(net20),
    .X(_0902_));
 sky130_fd_sc_hd__a221o_1 _1224_ (.A1(\a[27] ),
    .A2(net175),
    .B1(net158),
    .B2(\a[26] ),
    .C1(_0902_),
    .X(_0330_));
 sky130_fd_sc_hd__and2_1 _1225_ (.A(net201),
    .B(net19),
    .X(_0903_));
 sky130_fd_sc_hd__a221o_1 _1226_ (.A1(\a[26] ),
    .A2(net179),
    .B1(net162),
    .B2(\a[25] ),
    .C1(_0903_),
    .X(_0329_));
 sky130_fd_sc_hd__and2_1 _1227_ (.A(net201),
    .B(net18),
    .X(_0904_));
 sky130_fd_sc_hd__a221o_1 _1228_ (.A1(\a[25] ),
    .A2(net179),
    .B1(net162),
    .B2(\a[24] ),
    .C1(_0904_),
    .X(_0328_));
 sky130_fd_sc_hd__and2_1 _1229_ (.A(net201),
    .B(net17),
    .X(_0905_));
 sky130_fd_sc_hd__a221o_1 _1230_ (.A1(\a[24] ),
    .A2(net181),
    .B1(net164),
    .B2(\a[23] ),
    .C1(_0905_),
    .X(_0327_));
 sky130_fd_sc_hd__and2_1 _1231_ (.A(net201),
    .B(net16),
    .X(_0906_));
 sky130_fd_sc_hd__a221o_1 _1232_ (.A1(\a[23] ),
    .A2(net181),
    .B1(net164),
    .B2(\a[22] ),
    .C1(_0906_),
    .X(_0326_));
 sky130_fd_sc_hd__and2_1 _1233_ (.A(net201),
    .B(net15),
    .X(_0907_));
 sky130_fd_sc_hd__a221o_1 _1234_ (.A1(\a[22] ),
    .A2(net181),
    .B1(net164),
    .B2(\a[21] ),
    .C1(_0907_),
    .X(_0325_));
 sky130_fd_sc_hd__and2_1 _1235_ (.A(net201),
    .B(net14),
    .X(_0908_));
 sky130_fd_sc_hd__a221o_1 _1236_ (.A1(\a[21] ),
    .A2(net180),
    .B1(net163),
    .B2(\a[20] ),
    .C1(_0908_),
    .X(_0324_));
 sky130_fd_sc_hd__and2_1 _1237_ (.A(net201),
    .B(net13),
    .X(_0909_));
 sky130_fd_sc_hd__a221o_1 _1238_ (.A1(\a[20] ),
    .A2(net179),
    .B1(net162),
    .B2(\a[19] ),
    .C1(_0909_),
    .X(_0323_));
 sky130_fd_sc_hd__and2_1 _1239_ (.A(net200),
    .B(net11),
    .X(_0910_));
 sky130_fd_sc_hd__a221o_1 _1240_ (.A1(\a[19] ),
    .A2(net180),
    .B1(net163),
    .B2(\a[18] ),
    .C1(_0910_),
    .X(_0322_));
 sky130_fd_sc_hd__and2_1 _1241_ (.A(net200),
    .B(net10),
    .X(_0911_));
 sky130_fd_sc_hd__a221o_1 _1242_ (.A1(\a[18] ),
    .A2(net180),
    .B1(net163),
    .B2(\a[17] ),
    .C1(_0911_),
    .X(_0321_));
 sky130_fd_sc_hd__and2_1 _1243_ (.A(net200),
    .B(net9),
    .X(_0912_));
 sky130_fd_sc_hd__a221o_1 _1244_ (.A1(\a[17] ),
    .A2(net180),
    .B1(net163),
    .B2(\a[16] ),
    .C1(_0912_),
    .X(_0320_));
 sky130_fd_sc_hd__and2_1 _1245_ (.A(net200),
    .B(net8),
    .X(_0913_));
 sky130_fd_sc_hd__a221o_1 _1246_ (.A1(\a[16] ),
    .A2(net180),
    .B1(net163),
    .B2(\a[15] ),
    .C1(_0913_),
    .X(_0319_));
 sky130_fd_sc_hd__and2_1 _1247_ (.A(net200),
    .B(net7),
    .X(_0914_));
 sky130_fd_sc_hd__a221o_1 _1248_ (.A1(\a[15] ),
    .A2(net179),
    .B1(net162),
    .B2(\a[14] ),
    .C1(_0914_),
    .X(_0318_));
 sky130_fd_sc_hd__and2_1 _1249_ (.A(net201),
    .B(net6),
    .X(_0915_));
 sky130_fd_sc_hd__a221o_1 _1250_ (.A1(\a[14] ),
    .A2(net179),
    .B1(net162),
    .B2(\a[13] ),
    .C1(_0915_),
    .X(_0317_));
 sky130_fd_sc_hd__and2_1 _1251_ (.A(net200),
    .B(net5),
    .X(_0916_));
 sky130_fd_sc_hd__a221o_1 _1252_ (.A1(\a[13] ),
    .A2(net179),
    .B1(net162),
    .B2(\a[12] ),
    .C1(_0916_),
    .X(_0316_));
 sky130_fd_sc_hd__and2_1 _1253_ (.A(net200),
    .B(net4),
    .X(_0917_));
 sky130_fd_sc_hd__a221o_1 _1254_ (.A1(\a[12] ),
    .A2(net179),
    .B1(net162),
    .B2(\a[11] ),
    .C1(_0917_),
    .X(_0315_));
 sky130_fd_sc_hd__and2_1 _1255_ (.A(net200),
    .B(net3),
    .X(_0398_));
 sky130_fd_sc_hd__a221o_1 _1256_ (.A1(\a[11] ),
    .A2(net179),
    .B1(net162),
    .B2(\a[10] ),
    .C1(_0398_),
    .X(_0314_));
 sky130_fd_sc_hd__and2_1 _1257_ (.A(net200),
    .B(net2),
    .X(_0399_));
 sky130_fd_sc_hd__a221o_1 _1258_ (.A1(\a[10] ),
    .A2(net179),
    .B1(net162),
    .B2(\a[9] ),
    .C1(_0399_),
    .X(_0313_));
 sky130_fd_sc_hd__and2_1 _1259_ (.A(net200),
    .B(net32),
    .X(_0400_));
 sky130_fd_sc_hd__a221o_1 _1260_ (.A1(\a[9] ),
    .A2(net179),
    .B1(net162),
    .B2(\a[8] ),
    .C1(_0400_),
    .X(_0312_));
 sky130_fd_sc_hd__and2_1 _1261_ (.A(net198),
    .B(net31),
    .X(_0401_));
 sky130_fd_sc_hd__a221o_1 _1262_ (.A1(\a[8] ),
    .A2(net175),
    .B1(net158),
    .B2(\a[7] ),
    .C1(_0401_),
    .X(_0311_));
 sky130_fd_sc_hd__and2_1 _1263_ (.A(net198),
    .B(net30),
    .X(_0402_));
 sky130_fd_sc_hd__a221o_1 _1264_ (.A1(\a[7] ),
    .A2(net175),
    .B1(net158),
    .B2(\a[6] ),
    .C1(_0402_),
    .X(_0310_));
 sky130_fd_sc_hd__and2_1 _1265_ (.A(net196),
    .B(net29),
    .X(_0403_));
 sky130_fd_sc_hd__a221o_1 _1266_ (.A1(\a[6] ),
    .A2(net174),
    .B1(net157),
    .B2(\a[5] ),
    .C1(_0403_),
    .X(_0309_));
 sky130_fd_sc_hd__and2_1 _1267_ (.A(net196),
    .B(net28),
    .X(_0404_));
 sky130_fd_sc_hd__a221o_1 _1268_ (.A1(\a[5] ),
    .A2(net173),
    .B1(net156),
    .B2(\a[4] ),
    .C1(_0404_),
    .X(_0308_));
 sky130_fd_sc_hd__and2_1 _1269_ (.A(net196),
    .B(net27),
    .X(_0405_));
 sky130_fd_sc_hd__a221o_1 _1270_ (.A1(\a[4] ),
    .A2(net173),
    .B1(net156),
    .B2(\a[3] ),
    .C1(_0405_),
    .X(_0307_));
 sky130_fd_sc_hd__and2_1 _1271_ (.A(net196),
    .B(net26),
    .X(_0406_));
 sky130_fd_sc_hd__a221o_1 _1272_ (.A1(\a[3] ),
    .A2(net173),
    .B1(net156),
    .B2(\a[2] ),
    .C1(_0406_),
    .X(_0306_));
 sky130_fd_sc_hd__and2_1 _1273_ (.A(net199),
    .B(net23),
    .X(_0407_));
 sky130_fd_sc_hd__a221o_1 _1274_ (.A1(\a[2] ),
    .A2(net174),
    .B1(net157),
    .B2(\a[1] ),
    .C1(_0407_),
    .X(_0305_));
 sky130_fd_sc_hd__and2_1 _1275_ (.A(net196),
    .B(net12),
    .X(_0408_));
 sky130_fd_sc_hd__a221o_1 _1276_ (.A1(\a[1] ),
    .A2(net174),
    .B1(net157),
    .B2(\a[0] ),
    .C1(_0408_),
    .X(_0304_));
 sky130_fd_sc_hd__a22o_1 _1277_ (.A1(net202),
    .A2(net1),
    .B1(net176),
    .B2(\a[0] ),
    .X(_0303_));
 sky130_fd_sc_hd__a21oi_4 _1278_ (.A1(net57),
    .A2(net25),
    .B1(net168),
    .Y(_0409_));
 sky130_fd_sc_hd__a21o_1 _1279_ (.A1(\temp_product[63] ),
    .A2(net139),
    .B1(net149),
    .X(_0410_));
 sky130_fd_sc_hd__nand2_1 _1280_ (.A(net194),
    .B(\temp_product[62] ),
    .Y(_0411_));
 sky130_fd_sc_hd__xnor2_1 _1281_ (.A(net192),
    .B(\temp_product[56] ),
    .Y(_0412_));
 sky130_fd_sc_hd__nand2_1 _1282_ (.A(net194),
    .B(\temp_product[52] ),
    .Y(_0413_));
 sky130_fd_sc_hd__or2_1 _1283_ (.A(net193),
    .B(\temp_product[52] ),
    .X(_0414_));
 sky130_fd_sc_hd__and2_1 _1284_ (.A(_0413_),
    .B(_0414_),
    .X(_0415_));
 sky130_fd_sc_hd__and2_1 _1285_ (.A(net193),
    .B(\temp_product[54] ),
    .X(_0416_));
 sky130_fd_sc_hd__nor2_1 _1286_ (.A(net193),
    .B(\temp_product[54] ),
    .Y(_0417_));
 sky130_fd_sc_hd__nor2_1 _1287_ (.A(_0416_),
    .B(_0417_),
    .Y(_0418_));
 sky130_fd_sc_hd__xor2_1 _1288_ (.A(net193),
    .B(\temp_product[55] ),
    .X(_0419_));
 sky130_fd_sc_hd__xor2_1 _1289_ (.A(net194),
    .B(\temp_product[53] ),
    .X(_0420_));
 sky130_fd_sc_hd__and4_1 _1290_ (.A(_0415_),
    .B(_0418_),
    .C(_0419_),
    .D(_0420_),
    .X(_0421_));
 sky130_fd_sc_hd__nand2_1 _1291_ (.A(net195),
    .B(\temp_product[48] ),
    .Y(_0422_));
 sky130_fd_sc_hd__or2_1 _1292_ (.A(net195),
    .B(\temp_product[48] ),
    .X(_0423_));
 sky130_fd_sc_hd__nand2_1 _1293_ (.A(_0422_),
    .B(_0423_),
    .Y(_0424_));
 sky130_fd_sc_hd__xor2_1 _1294_ (.A(net195),
    .B(\temp_product[51] ),
    .X(_0425_));
 sky130_fd_sc_hd__nand2_1 _1295_ (.A(net195),
    .B(\temp_product[50] ),
    .Y(_0426_));
 sky130_fd_sc_hd__or2_1 _1296_ (.A(net195),
    .B(\temp_product[50] ),
    .X(_0427_));
 sky130_fd_sc_hd__and2_1 _1297_ (.A(_0426_),
    .B(_0427_),
    .X(_0428_));
 sky130_fd_sc_hd__xor2_2 _1298_ (.A(net195),
    .B(\temp_product[49] ),
    .X(_0429_));
 sky130_fd_sc_hd__nand4b_1 _1299_ (.A_N(_0424_),
    .B(_0425_),
    .C(_0428_),
    .D(_0429_),
    .Y(_0430_));
 sky130_fd_sc_hd__or4_1 _1300_ (.A(_0679_),
    .B(_0682_),
    .C(_0688_),
    .D(_0801_),
    .X(_0431_));
 sky130_fd_sc_hd__nor3_1 _1301_ (.A(_0694_),
    .B(_0696_),
    .C(_0431_),
    .Y(_0432_));
 sky130_fd_sc_hd__and3_1 _1302_ (.A(_0700_),
    .B(_0808_),
    .C(_0432_),
    .X(_0433_));
 sky130_fd_sc_hd__and2_1 _1303_ (.A(_0789_),
    .B(_0433_),
    .X(_0434_));
 sky130_fd_sc_hd__o211a_1 _1304_ (.A1(\temp_product[25] ),
    .A2(\a[25] ),
    .B1(_0698_),
    .C1(_0432_),
    .X(_0435_));
 sky130_fd_sc_hd__or4_1 _1305_ (.A(_0679_),
    .B(_0682_),
    .C(_0683_),
    .D(_0686_),
    .X(_0436_));
 sky130_fd_sc_hd__and3_1 _1306_ (.A(\temp_product[30] ),
    .B(\a[30] ),
    .C(_0678_),
    .X(_0437_));
 sky130_fd_sc_hd__o21ai_1 _1307_ (.A1(_0693_),
    .A2(_0431_),
    .B1(_0436_),
    .Y(_0438_));
 sky130_fd_sc_hd__or4b_1 _1308_ (.A(_0435_),
    .B(_0438_),
    .C(_0437_),
    .D_N(_0677_),
    .X(_0439_));
 sky130_fd_sc_hd__a21o_1 _1309_ (.A1(_0730_),
    .A2(_0433_),
    .B1(_0439_),
    .X(_0440_));
 sky130_fd_sc_hd__a21o_2 _1310_ (.A1(_0786_),
    .A2(_0434_),
    .B1(_0440_),
    .X(_0441_));
 sky130_fd_sc_hd__xor2_1 _1311_ (.A(net189),
    .B(\temp_product[35] ),
    .X(_0442_));
 sky130_fd_sc_hd__nand2_1 _1312_ (.A(net189),
    .B(\temp_product[32] ),
    .Y(_0443_));
 sky130_fd_sc_hd__or2_1 _1313_ (.A(net189),
    .B(\temp_product[32] ),
    .X(_0444_));
 sky130_fd_sc_hd__and2_1 _1314_ (.A(_0443_),
    .B(_0444_),
    .X(_0445_));
 sky130_fd_sc_hd__nand2_1 _1315_ (.A(net189),
    .B(\temp_product[34] ),
    .Y(_0446_));
 sky130_fd_sc_hd__or2_1 _1316_ (.A(net189),
    .B(\temp_product[34] ),
    .X(_0447_));
 sky130_fd_sc_hd__nand2_1 _1317_ (.A(_0446_),
    .B(_0447_),
    .Y(_0448_));
 sky130_fd_sc_hd__xor2_2 _1318_ (.A(net189),
    .B(\temp_product[33] ),
    .X(_0449_));
 sky130_fd_sc_hd__and3_1 _1319_ (.A(_0442_),
    .B(_0446_),
    .C(_0447_),
    .X(_0450_));
 sky130_fd_sc_hd__nand2_1 _1320_ (.A(net187),
    .B(\temp_product[38] ),
    .Y(_0451_));
 sky130_fd_sc_hd__or2_1 _1321_ (.A(net187),
    .B(\temp_product[38] ),
    .X(_0452_));
 sky130_fd_sc_hd__nand2_1 _1322_ (.A(_0451_),
    .B(_0452_),
    .Y(_0453_));
 sky130_fd_sc_hd__xor2_1 _1323_ (.A(net187),
    .B(\temp_product[39] ),
    .X(_0454_));
 sky130_fd_sc_hd__nand2_1 _1324_ (.A(net187),
    .B(\temp_product[36] ),
    .Y(_0455_));
 sky130_fd_sc_hd__or2_1 _1325_ (.A(net187),
    .B(\temp_product[36] ),
    .X(_0456_));
 sky130_fd_sc_hd__nand2_1 _1326_ (.A(_0455_),
    .B(_0456_),
    .Y(_0457_));
 sky130_fd_sc_hd__inv_2 _1327_ (.A(_0457_),
    .Y(_0458_));
 sky130_fd_sc_hd__nand2_1 _1328_ (.A(net187),
    .B(\temp_product[37] ),
    .Y(_0459_));
 sky130_fd_sc_hd__or2_1 _1329_ (.A(net191),
    .B(\temp_product[37] ),
    .X(_0460_));
 sky130_fd_sc_hd__and2_1 _1330_ (.A(_0459_),
    .B(_0460_),
    .X(_0461_));
 sky130_fd_sc_hd__and4b_1 _1331_ (.A_N(_0453_),
    .B(_0454_),
    .C(_0458_),
    .D(_0461_),
    .X(_0462_));
 sky130_fd_sc_hd__and4_1 _1332_ (.A(_0445_),
    .B(_0449_),
    .C(_0450_),
    .D(_0462_),
    .X(_0463_));
 sky130_fd_sc_hd__nand2_1 _1333_ (.A(_0441_),
    .B(_0463_),
    .Y(_0464_));
 sky130_fd_sc_hd__nand2_1 _1334_ (.A(net188),
    .B(\temp_product[43] ),
    .Y(_0465_));
 sky130_fd_sc_hd__or2_1 _1335_ (.A(net188),
    .B(\temp_product[43] ),
    .X(_0466_));
 sky130_fd_sc_hd__and2_1 _1336_ (.A(_0465_),
    .B(_0466_),
    .X(_0467_));
 sky130_fd_sc_hd__nand2_1 _1337_ (.A(net188),
    .B(\temp_product[42] ),
    .Y(_0468_));
 sky130_fd_sc_hd__or2_1 _1338_ (.A(net188),
    .B(\temp_product[42] ),
    .X(_0469_));
 sky130_fd_sc_hd__nand2_1 _1339_ (.A(_0468_),
    .B(_0469_),
    .Y(_0470_));
 sky130_fd_sc_hd__xor2_1 _1340_ (.A(net188),
    .B(\temp_product[41] ),
    .X(_0471_));
 sky130_fd_sc_hd__and4_1 _1341_ (.A(_0467_),
    .B(_0468_),
    .C(_0469_),
    .D(_0471_),
    .X(_0472_));
 sky130_fd_sc_hd__xor2_1 _1342_ (.A(net190),
    .B(\temp_product[45] ),
    .X(_0473_));
 sky130_fd_sc_hd__inv_2 _1343_ (.A(_0473_),
    .Y(_0474_));
 sky130_fd_sc_hd__xnor2_1 _1344_ (.A(net187),
    .B(\temp_product[40] ),
    .Y(_0475_));
 sky130_fd_sc_hd__xor2_1 _1345_ (.A(net190),
    .B(\temp_product[47] ),
    .X(_0476_));
 sky130_fd_sc_hd__nand2_1 _1346_ (.A(net189),
    .B(\temp_product[46] ),
    .Y(_0477_));
 sky130_fd_sc_hd__or2_1 _1347_ (.A(net190),
    .B(\temp_product[46] ),
    .X(_0478_));
 sky130_fd_sc_hd__nand2_1 _1348_ (.A(_0477_),
    .B(_0478_),
    .Y(_0479_));
 sky130_fd_sc_hd__nand2_1 _1349_ (.A(net190),
    .B(\temp_product[44] ),
    .Y(_0480_));
 sky130_fd_sc_hd__or2_1 _1350_ (.A(net187),
    .B(\temp_product[44] ),
    .X(_0481_));
 sky130_fd_sc_hd__nand2_1 _1351_ (.A(_0480_),
    .B(_0481_),
    .Y(_0482_));
 sky130_fd_sc_hd__nor2_1 _1352_ (.A(_0475_),
    .B(_0482_),
    .Y(_0483_));
 sky130_fd_sc_hd__nor2_1 _1353_ (.A(_0474_),
    .B(_0479_),
    .Y(_0484_));
 sky130_fd_sc_hd__and4_1 _1354_ (.A(_0472_),
    .B(_0476_),
    .C(_0483_),
    .D(_0484_),
    .X(_0485_));
 sky130_fd_sc_hd__o21a_1 _1355_ (.A1(\temp_product[33] ),
    .A2(\temp_product[32] ),
    .B1(net189),
    .X(_0486_));
 sky130_fd_sc_hd__o41a_1 _1356_ (.A1(\temp_product[35] ),
    .A2(\temp_product[34] ),
    .A3(\temp_product[33] ),
    .A4(\temp_product[32] ),
    .B1(net189),
    .X(_0487_));
 sky130_fd_sc_hd__o41a_1 _1357_ (.A1(\temp_product[39] ),
    .A2(\temp_product[38] ),
    .A3(\temp_product[37] ),
    .A4(\temp_product[36] ),
    .B1(net187),
    .X(_0488_));
 sky130_fd_sc_hd__nor2_1 _1358_ (.A(_0487_),
    .B(_0488_),
    .Y(_0489_));
 sky130_fd_sc_hd__o21ai_1 _1359_ (.A1(\temp_product[41] ),
    .A2(\temp_product[40] ),
    .B1(net187),
    .Y(_0490_));
 sky130_fd_sc_hd__and3_1 _1360_ (.A(_0465_),
    .B(_0468_),
    .C(_0490_),
    .X(_0491_));
 sky130_fd_sc_hd__o21ai_2 _1361_ (.A1(\temp_product[45] ),
    .A2(\temp_product[44] ),
    .B1(net190),
    .Y(_0492_));
 sky130_fd_sc_hd__o21ai_1 _1362_ (.A1(\temp_product[47] ),
    .A2(\temp_product[46] ),
    .B1(net189),
    .Y(_0493_));
 sky130_fd_sc_hd__nand4_2 _1363_ (.A(_0489_),
    .B(_0491_),
    .C(_0492_),
    .D(_0493_),
    .Y(_0494_));
 sky130_fd_sc_hd__a31oi_4 _1364_ (.A1(_0441_),
    .A2(_0463_),
    .A3(_0485_),
    .B1(_0494_),
    .Y(_0495_));
 sky130_fd_sc_hd__nor2_1 _1365_ (.A(_0430_),
    .B(_0495_),
    .Y(_0496_));
 sky130_fd_sc_hd__or3b_1 _1366_ (.A(_0495_),
    .B(_0430_),
    .C_N(_0421_),
    .X(_0497_));
 sky130_fd_sc_hd__o21a_1 _1367_ (.A1(\temp_product[49] ),
    .A2(\temp_product[48] ),
    .B1(net195),
    .X(_0498_));
 sky130_fd_sc_hd__o41a_1 _1368_ (.A1(\temp_product[51] ),
    .A2(\temp_product[50] ),
    .A3(\temp_product[49] ),
    .A4(\temp_product[48] ),
    .B1(net195),
    .X(_0499_));
 sky130_fd_sc_hd__o21a_1 _1369_ (.A1(\temp_product[53] ),
    .A2(\temp_product[52] ),
    .B1(net193),
    .X(_0500_));
 sky130_fd_sc_hd__a2111oi_1 _1370_ (.A1(net193),
    .A2(\temp_product[55] ),
    .B1(_0416_),
    .C1(_0499_),
    .D1(_0500_),
    .Y(_0501_));
 sky130_fd_sc_hd__nand2_1 _1371_ (.A(_0497_),
    .B(_0501_),
    .Y(_0502_));
 sky130_fd_sc_hd__a21oi_1 _1372_ (.A1(_0497_),
    .A2(net186),
    .B1(_0412_),
    .Y(_0503_));
 sky130_fd_sc_hd__nand2_1 _1373_ (.A(net192),
    .B(\temp_product[58] ),
    .Y(_0504_));
 sky130_fd_sc_hd__or2_1 _1374_ (.A(net192),
    .B(\temp_product[58] ),
    .X(_0505_));
 sky130_fd_sc_hd__nand2_1 _1375_ (.A(_0504_),
    .B(_0505_),
    .Y(_0506_));
 sky130_fd_sc_hd__xor2_1 _1376_ (.A(net193),
    .B(\temp_product[59] ),
    .X(_0507_));
 sky130_fd_sc_hd__xor2_1 _1377_ (.A(net192),
    .B(\temp_product[57] ),
    .X(_0508_));
 sky130_fd_sc_hd__and4_1 _1378_ (.A(_0504_),
    .B(_0505_),
    .C(_0507_),
    .D(_0508_),
    .X(_0509_));
 sky130_fd_sc_hd__nand2_1 _1379_ (.A(_0503_),
    .B(_0508_),
    .Y(_0510_));
 sky130_fd_sc_hd__o21ai_1 _1380_ (.A1(\temp_product[57] ),
    .A2(\temp_product[56] ),
    .B1(net192),
    .Y(_0511_));
 sky130_fd_sc_hd__o41a_1 _1381_ (.A1(\temp_product[59] ),
    .A2(\temp_product[58] ),
    .A3(\temp_product[57] ),
    .A4(\temp_product[56] ),
    .B1(net192),
    .X(_0512_));
 sky130_fd_sc_hd__a21o_1 _1382_ (.A1(_0503_),
    .A2(_0509_),
    .B1(_0512_),
    .X(_0513_));
 sky130_fd_sc_hd__and2_1 _1383_ (.A(net192),
    .B(\temp_product[60] ),
    .X(_0514_));
 sky130_fd_sc_hd__nor2_1 _1384_ (.A(net192),
    .B(\temp_product[60] ),
    .Y(_0515_));
 sky130_fd_sc_hd__nor2_1 _1385_ (.A(_0514_),
    .B(_0515_),
    .Y(_0516_));
 sky130_fd_sc_hd__xor2_1 _1386_ (.A(net194),
    .B(\temp_product[61] ),
    .X(_0517_));
 sky130_fd_sc_hd__o21a_1 _1387_ (.A1(\temp_product[61] ),
    .A2(\temp_product[60] ),
    .B1(net192),
    .X(_0518_));
 sky130_fd_sc_hd__a31o_1 _1388_ (.A1(_0513_),
    .A2(_0516_),
    .A3(_0517_),
    .B1(_0518_),
    .X(_0519_));
 sky130_fd_sc_hd__or2_1 _1389_ (.A(net194),
    .B(\temp_product[62] ),
    .X(_0520_));
 sky130_fd_sc_hd__and3_1 _1390_ (.A(_0411_),
    .B(_0519_),
    .C(_0520_),
    .X(_0521_));
 sky130_fd_sc_hd__a21boi_1 _1391_ (.A1(_0519_),
    .A2(_0520_),
    .B1_N(_0411_),
    .Y(_0522_));
 sky130_fd_sc_hd__or2_1 _1392_ (.A(net194),
    .B(\temp_product[63] ),
    .X(_0523_));
 sky130_fd_sc_hd__nand2_1 _1393_ (.A(net194),
    .B(\temp_product[63] ),
    .Y(_0524_));
 sky130_fd_sc_hd__a21oi_1 _1394_ (.A1(_0523_),
    .A2(_0524_),
    .B1(_0522_),
    .Y(_0525_));
 sky130_fd_sc_hd__a31o_1 _1395_ (.A1(_0522_),
    .A2(_0523_),
    .A3(_0524_),
    .B1(_0669_),
    .X(_0526_));
 sky130_fd_sc_hd__or2_1 _1396_ (.A(_0525_),
    .B(_0526_),
    .X(_0527_));
 sky130_fd_sc_hd__a22o_1 _1397_ (.A1(\temp_product[63] ),
    .A2(net154),
    .B1(_0410_),
    .B2(_0527_),
    .X(_0302_));
 sky130_fd_sc_hd__a21oi_1 _1398_ (.A1(_0411_),
    .A2(_0520_),
    .B1(_0519_),
    .Y(_0528_));
 sky130_fd_sc_hd__o21ai_1 _1399_ (.A1(_0521_),
    .A2(_0528_),
    .B1(net182),
    .Y(_0529_));
 sky130_fd_sc_hd__a21o_1 _1400_ (.A1(\temp_product[62] ),
    .A2(net139),
    .B1(net149),
    .X(_0530_));
 sky130_fd_sc_hd__a22o_1 _1401_ (.A1(\temp_product[62] ),
    .A2(net154),
    .B1(_0529_),
    .B2(_0530_),
    .X(_0301_));
 sky130_fd_sc_hd__a21o_1 _1402_ (.A1(\temp_product[61] ),
    .A2(net138),
    .B1(net149),
    .X(_0531_));
 sky130_fd_sc_hd__nand2_1 _1403_ (.A(_0513_),
    .B(_0516_),
    .Y(_0532_));
 sky130_fd_sc_hd__a21oi_1 _1404_ (.A1(_0513_),
    .A2(_0516_),
    .B1(_0514_),
    .Y(_0533_));
 sky130_fd_sc_hd__o21ai_1 _1405_ (.A1(_0517_),
    .A2(_0533_),
    .B1(net182),
    .Y(_0534_));
 sky130_fd_sc_hd__a21o_1 _1406_ (.A1(_0517_),
    .A2(_0533_),
    .B1(_0534_),
    .X(_0535_));
 sky130_fd_sc_hd__a22o_1 _1407_ (.A1(\temp_product[61] ),
    .A2(net154),
    .B1(_0531_),
    .B2(_0535_),
    .X(_0300_));
 sky130_fd_sc_hd__or2_1 _1408_ (.A(_0513_),
    .B(_0516_),
    .X(_0536_));
 sky130_fd_sc_hd__a21o_1 _1409_ (.A1(_0532_),
    .A2(_0536_),
    .B1(net185),
    .X(_0537_));
 sky130_fd_sc_hd__a21o_1 _1410_ (.A1(\temp_product[60] ),
    .A2(net142),
    .B1(net150),
    .X(_0538_));
 sky130_fd_sc_hd__a22o_1 _1411_ (.A1(\temp_product[60] ),
    .A2(net155),
    .B1(_0537_),
    .B2(_0538_),
    .X(_0299_));
 sky130_fd_sc_hd__a21o_1 _1412_ (.A1(\temp_product[59] ),
    .A2(net142),
    .B1(net150),
    .X(_0539_));
 sky130_fd_sc_hd__a21o_1 _1413_ (.A1(_0510_),
    .A2(_0511_),
    .B1(_0506_),
    .X(_0540_));
 sky130_fd_sc_hd__and3_1 _1414_ (.A(_0504_),
    .B(_0507_),
    .C(_0540_),
    .X(_0541_));
 sky130_fd_sc_hd__a21oi_1 _1415_ (.A1(_0504_),
    .A2(_0540_),
    .B1(_0507_),
    .Y(_0542_));
 sky130_fd_sc_hd__or3_1 _1416_ (.A(net185),
    .B(_0541_),
    .C(_0542_),
    .X(_0543_));
 sky130_fd_sc_hd__a22o_1 _1417_ (.A1(\temp_product[59] ),
    .A2(net154),
    .B1(_0539_),
    .B2(_0543_),
    .X(_0298_));
 sky130_fd_sc_hd__nand3_1 _1418_ (.A(_0506_),
    .B(_0510_),
    .C(_0511_),
    .Y(_0544_));
 sky130_fd_sc_hd__a21o_1 _1419_ (.A1(_0540_),
    .A2(_0544_),
    .B1(net185),
    .X(_0545_));
 sky130_fd_sc_hd__a21o_1 _1420_ (.A1(\temp_product[58] ),
    .A2(net142),
    .B1(net149),
    .X(_0546_));
 sky130_fd_sc_hd__a22o_1 _1421_ (.A1(\temp_product[58] ),
    .A2(net154),
    .B1(_0545_),
    .B2(_0546_),
    .X(_0297_));
 sky130_fd_sc_hd__a21o_1 _1422_ (.A1(\temp_product[57] ),
    .A2(net142),
    .B1(net149),
    .X(_0547_));
 sky130_fd_sc_hd__a21oi_1 _1423_ (.A1(net192),
    .A2(\temp_product[56] ),
    .B1(_0503_),
    .Y(_0548_));
 sky130_fd_sc_hd__a21oi_1 _1424_ (.A1(_0508_),
    .A2(_0548_),
    .B1(net185),
    .Y(_0549_));
 sky130_fd_sc_hd__o21ai_1 _1425_ (.A1(_0508_),
    .A2(_0548_),
    .B1(_0549_),
    .Y(_0550_));
 sky130_fd_sc_hd__a22o_1 _1426_ (.A1(\temp_product[57] ),
    .A2(net154),
    .B1(_0547_),
    .B2(_0550_),
    .X(_0296_));
 sky130_fd_sc_hd__xor2_1 _1427_ (.A(_0412_),
    .B(_0502_),
    .X(_0551_));
 sky130_fd_sc_hd__nand2_1 _1428_ (.A(net182),
    .B(_0551_),
    .Y(_0552_));
 sky130_fd_sc_hd__a21o_1 _1429_ (.A1(\temp_product[56] ),
    .A2(net142),
    .B1(net149),
    .X(_0553_));
 sky130_fd_sc_hd__a22o_1 _1430_ (.A1(\temp_product[56] ),
    .A2(net154),
    .B1(_0552_),
    .B2(_0553_),
    .X(_0295_));
 sky130_fd_sc_hd__a21o_1 _1431_ (.A1(\temp_product[55] ),
    .A2(net141),
    .B1(net149),
    .X(_0554_));
 sky130_fd_sc_hd__o21ai_2 _1432_ (.A1(_0496_),
    .A2(_0499_),
    .B1(_0415_),
    .Y(_0555_));
 sky130_fd_sc_hd__inv_2 _1433_ (.A(_0555_),
    .Y(_0556_));
 sky130_fd_sc_hd__a21o_1 _1434_ (.A1(_0420_),
    .A2(_0556_),
    .B1(_0500_),
    .X(_0557_));
 sky130_fd_sc_hd__a21o_1 _1435_ (.A1(_0418_),
    .A2(_0557_),
    .B1(_0416_),
    .X(_0558_));
 sky130_fd_sc_hd__xnor2_1 _1436_ (.A(_0419_),
    .B(_0558_),
    .Y(_0559_));
 sky130_fd_sc_hd__nand2_1 _1437_ (.A(net182),
    .B(_0559_),
    .Y(_0560_));
 sky130_fd_sc_hd__a22o_1 _1438_ (.A1(\temp_product[55] ),
    .A2(net154),
    .B1(_0554_),
    .B2(_0560_),
    .X(_0294_));
 sky130_fd_sc_hd__xnor2_1 _1439_ (.A(_0418_),
    .B(_0557_),
    .Y(_0561_));
 sky130_fd_sc_hd__nand2_1 _1440_ (.A(net182),
    .B(_0561_),
    .Y(_0562_));
 sky130_fd_sc_hd__a21o_1 _1441_ (.A1(\temp_product[54] ),
    .A2(net141),
    .B1(net150),
    .X(_0563_));
 sky130_fd_sc_hd__a22o_1 _1442_ (.A1(\temp_product[54] ),
    .A2(net155),
    .B1(_0562_),
    .B2(_0563_),
    .X(_0293_));
 sky130_fd_sc_hd__a21o_1 _1443_ (.A1(\temp_product[53] ),
    .A2(net142),
    .B1(net149),
    .X(_0564_));
 sky130_fd_sc_hd__a21oi_1 _1444_ (.A1(_0413_),
    .A2(_0555_),
    .B1(_0420_),
    .Y(_0565_));
 sky130_fd_sc_hd__a31o_1 _1445_ (.A1(_0413_),
    .A2(_0420_),
    .A3(_0555_),
    .B1(net185),
    .X(_0566_));
 sky130_fd_sc_hd__or2_1 _1446_ (.A(_0565_),
    .B(_0566_),
    .X(_0567_));
 sky130_fd_sc_hd__a22o_1 _1447_ (.A1(\temp_product[53] ),
    .A2(net154),
    .B1(_0564_),
    .B2(_0567_),
    .X(_0292_));
 sky130_fd_sc_hd__or3_1 _1448_ (.A(_0415_),
    .B(_0496_),
    .C(_0499_),
    .X(_0568_));
 sky130_fd_sc_hd__a21o_1 _1449_ (.A1(_0555_),
    .A2(_0568_),
    .B1(net185),
    .X(_0569_));
 sky130_fd_sc_hd__a21o_1 _1450_ (.A1(\temp_product[52] ),
    .A2(net140),
    .B1(net150),
    .X(_0570_));
 sky130_fd_sc_hd__a22o_1 _1451_ (.A1(\temp_product[52] ),
    .A2(net155),
    .B1(_0569_),
    .B2(_0570_),
    .X(_0291_));
 sky130_fd_sc_hd__a21o_1 _1452_ (.A1(\temp_product[51] ),
    .A2(net141),
    .B1(net150),
    .X(_0571_));
 sky130_fd_sc_hd__or2_1 _1453_ (.A(_0424_),
    .B(_0495_),
    .X(_0572_));
 sky130_fd_sc_hd__inv_2 _1454_ (.A(_0572_),
    .Y(_0573_));
 sky130_fd_sc_hd__a21o_1 _1455_ (.A1(_0429_),
    .A2(_0573_),
    .B1(_0498_),
    .X(_0574_));
 sky130_fd_sc_hd__a21bo_1 _1456_ (.A1(_0428_),
    .A2(_0574_),
    .B1_N(_0426_),
    .X(_0575_));
 sky130_fd_sc_hd__xnor2_1 _1457_ (.A(_0425_),
    .B(_0575_),
    .Y(_0576_));
 sky130_fd_sc_hd__nand2_1 _1458_ (.A(_0670_),
    .B(_0576_),
    .Y(_0577_));
 sky130_fd_sc_hd__a22o_1 _1459_ (.A1(\temp_product[51] ),
    .A2(net155),
    .B1(_0571_),
    .B2(_0577_),
    .X(_0290_));
 sky130_fd_sc_hd__xnor2_1 _1460_ (.A(_0428_),
    .B(_0574_),
    .Y(_0578_));
 sky130_fd_sc_hd__nand2_1 _1461_ (.A(net182),
    .B(_0578_),
    .Y(_0579_));
 sky130_fd_sc_hd__a21o_1 _1462_ (.A1(\temp_product[50] ),
    .A2(net141),
    .B1(net150),
    .X(_0580_));
 sky130_fd_sc_hd__a22o_1 _1463_ (.A1(\temp_product[50] ),
    .A2(net155),
    .B1(_0579_),
    .B2(_0580_),
    .X(_0289_));
 sky130_fd_sc_hd__a21o_1 _1464_ (.A1(\temp_product[49] ),
    .A2(net140),
    .B1(net150),
    .X(_0581_));
 sky130_fd_sc_hd__a21o_1 _1465_ (.A1(_0422_),
    .A2(_0572_),
    .B1(_0429_),
    .X(_0582_));
 sky130_fd_sc_hd__nand2_1 _1466_ (.A(net182),
    .B(_0582_),
    .Y(_0583_));
 sky130_fd_sc_hd__a31o_1 _1467_ (.A1(_0422_),
    .A2(_0429_),
    .A3(_0572_),
    .B1(_0583_),
    .X(_0584_));
 sky130_fd_sc_hd__a22o_1 _1468_ (.A1(\temp_product[49] ),
    .A2(net155),
    .B1(_0581_),
    .B2(_0584_),
    .X(_0288_));
 sky130_fd_sc_hd__nand2_1 _1469_ (.A(_0424_),
    .B(_0495_),
    .Y(_0585_));
 sky130_fd_sc_hd__a21o_1 _1470_ (.A1(_0572_),
    .A2(_0585_),
    .B1(net185),
    .X(_0586_));
 sky130_fd_sc_hd__a21o_1 _1471_ (.A1(\temp_product[48] ),
    .A2(net140),
    .B1(net150),
    .X(_0587_));
 sky130_fd_sc_hd__a22o_1 _1472_ (.A1(\temp_product[48] ),
    .A2(net155),
    .B1(_0586_),
    .B2(_0587_),
    .X(_0287_));
 sky130_fd_sc_hd__a21o_1 _1473_ (.A1(\temp_product[47] ),
    .A2(net138),
    .B1(net149),
    .X(_0588_));
 sky130_fd_sc_hd__nand2_1 _1474_ (.A(_0464_),
    .B(_0489_),
    .Y(_0589_));
 sky130_fd_sc_hd__a21oi_1 _1475_ (.A1(_0464_),
    .A2(_0489_),
    .B1(_0475_),
    .Y(_0590_));
 sky130_fd_sc_hd__nand2_1 _1476_ (.A(_0472_),
    .B(_0590_),
    .Y(_0591_));
 sky130_fd_sc_hd__a21o_1 _1477_ (.A1(_0491_),
    .A2(_0591_),
    .B1(_0482_),
    .X(_0592_));
 sky130_fd_sc_hd__or2_1 _1478_ (.A(_0474_),
    .B(_0592_),
    .X(_0593_));
 sky130_fd_sc_hd__a21o_1 _1479_ (.A1(_0492_),
    .A2(_0593_),
    .B1(_0479_),
    .X(_0594_));
 sky130_fd_sc_hd__a21oi_1 _1480_ (.A1(_0477_),
    .A2(_0594_),
    .B1(_0476_),
    .Y(_0595_));
 sky130_fd_sc_hd__a31o_1 _1481_ (.A1(_0476_),
    .A2(_0477_),
    .A3(_0594_),
    .B1(net184),
    .X(_0596_));
 sky130_fd_sc_hd__or2_1 _1482_ (.A(_0595_),
    .B(_0596_),
    .X(_0597_));
 sky130_fd_sc_hd__a22o_1 _1483_ (.A1(\temp_product[47] ),
    .A2(net153),
    .B1(_0588_),
    .B2(_0597_),
    .X(_0286_));
 sky130_fd_sc_hd__nand3_1 _1484_ (.A(_0479_),
    .B(_0492_),
    .C(_0593_),
    .Y(_0598_));
 sky130_fd_sc_hd__and2_1 _1485_ (.A(_0594_),
    .B(_0598_),
    .X(_0599_));
 sky130_fd_sc_hd__and2_1 _1486_ (.A(\temp_product[46] ),
    .B(net138),
    .X(_0600_));
 sky130_fd_sc_hd__o22a_1 _1487_ (.A1(net184),
    .A2(_0599_),
    .B1(_0600_),
    .B2(net148),
    .X(_0601_));
 sky130_fd_sc_hd__a21o_1 _1488_ (.A1(\temp_product[46] ),
    .A2(net153),
    .B1(_0601_),
    .X(_0285_));
 sky130_fd_sc_hd__a21o_1 _1489_ (.A1(\temp_product[45] ),
    .A2(_0409_),
    .B1(net148),
    .X(_0602_));
 sky130_fd_sc_hd__and3_1 _1490_ (.A(_0473_),
    .B(_0480_),
    .C(_0592_),
    .X(_0603_));
 sky130_fd_sc_hd__a21oi_1 _1491_ (.A1(_0480_),
    .A2(_0592_),
    .B1(_0473_),
    .Y(_0604_));
 sky130_fd_sc_hd__or3_1 _1492_ (.A(net184),
    .B(_0603_),
    .C(_0604_),
    .X(_0605_));
 sky130_fd_sc_hd__a22o_1 _1493_ (.A1(\temp_product[45] ),
    .A2(net153),
    .B1(_0602_),
    .B2(_0605_),
    .X(_0284_));
 sky130_fd_sc_hd__nand3_1 _1494_ (.A(_0482_),
    .B(_0491_),
    .C(_0591_),
    .Y(_0606_));
 sky130_fd_sc_hd__a21o_1 _1495_ (.A1(_0592_),
    .A2(_0606_),
    .B1(net184),
    .X(_0607_));
 sky130_fd_sc_hd__a21o_1 _1496_ (.A1(\temp_product[44] ),
    .A2(net137),
    .B1(net148),
    .X(_0608_));
 sky130_fd_sc_hd__a22o_1 _1497_ (.A1(\temp_product[44] ),
    .A2(net153),
    .B1(_0607_),
    .B2(_0608_),
    .X(_0283_));
 sky130_fd_sc_hd__a21o_1 _1498_ (.A1(\temp_product[43] ),
    .A2(net136),
    .B1(net151),
    .X(_0609_));
 sky130_fd_sc_hd__nand2_1 _1499_ (.A(_0471_),
    .B(_0590_),
    .Y(_0610_));
 sky130_fd_sc_hd__a21o_1 _1500_ (.A1(_0490_),
    .A2(_0610_),
    .B1(_0470_),
    .X(_0611_));
 sky130_fd_sc_hd__a21oi_1 _1501_ (.A1(_0468_),
    .A2(_0611_),
    .B1(_0467_),
    .Y(_0612_));
 sky130_fd_sc_hd__a31o_1 _1502_ (.A1(_0467_),
    .A2(_0468_),
    .A3(_0611_),
    .B1(net184),
    .X(_0613_));
 sky130_fd_sc_hd__or2_1 _1503_ (.A(_0612_),
    .B(_0613_),
    .X(_0614_));
 sky130_fd_sc_hd__a22o_1 _1504_ (.A1(\temp_product[43] ),
    .A2(net153),
    .B1(_0609_),
    .B2(_0614_),
    .X(_0282_));
 sky130_fd_sc_hd__nand3_1 _1505_ (.A(_0470_),
    .B(_0490_),
    .C(_0610_),
    .Y(_0615_));
 sky130_fd_sc_hd__a21o_1 _1506_ (.A1(_0611_),
    .A2(_0615_),
    .B1(net183),
    .X(_0616_));
 sky130_fd_sc_hd__a21o_1 _1507_ (.A1(\temp_product[42] ),
    .A2(net137),
    .B1(net151),
    .X(_0617_));
 sky130_fd_sc_hd__a22o_1 _1508_ (.A1(\temp_product[42] ),
    .A2(net152),
    .B1(_0616_),
    .B2(_0617_),
    .X(_0281_));
 sky130_fd_sc_hd__a21o_1 _1509_ (.A1(\temp_product[41] ),
    .A2(net136),
    .B1(net151),
    .X(_0618_));
 sky130_fd_sc_hd__a21oi_1 _1510_ (.A1(net188),
    .A2(\temp_product[40] ),
    .B1(_0590_),
    .Y(_0619_));
 sky130_fd_sc_hd__o21ai_1 _1511_ (.A1(_0471_),
    .A2(_0619_),
    .B1(net182),
    .Y(_0620_));
 sky130_fd_sc_hd__a21o_1 _1512_ (.A1(_0471_),
    .A2(_0619_),
    .B1(_0620_),
    .X(_0621_));
 sky130_fd_sc_hd__a22o_1 _1513_ (.A1(\temp_product[41] ),
    .A2(net152),
    .B1(_0618_),
    .B2(_0621_),
    .X(_0280_));
 sky130_fd_sc_hd__xnor2_1 _1514_ (.A(_0475_),
    .B(_0589_),
    .Y(_0622_));
 sky130_fd_sc_hd__or2_1 _1515_ (.A(net183),
    .B(_0622_),
    .X(_0623_));
 sky130_fd_sc_hd__a21o_1 _1516_ (.A1(\temp_product[40] ),
    .A2(net137),
    .B1(net148),
    .X(_0624_));
 sky130_fd_sc_hd__a22o_1 _1517_ (.A1(\temp_product[40] ),
    .A2(net152),
    .B1(_0623_),
    .B2(_0624_),
    .X(_0279_));
 sky130_fd_sc_hd__a21o_1 _1518_ (.A1(\temp_product[39] ),
    .A2(net137),
    .B1(net148),
    .X(_0625_));
 sky130_fd_sc_hd__nand2_1 _1519_ (.A(_0441_),
    .B(_0445_),
    .Y(_0626_));
 sky130_fd_sc_hd__inv_2 _1520_ (.A(_0626_),
    .Y(_0627_));
 sky130_fd_sc_hd__a31oi_2 _1521_ (.A1(_0449_),
    .A2(_0450_),
    .A3(_0627_),
    .B1(_0487_),
    .Y(_0628_));
 sky130_fd_sc_hd__or2_1 _1522_ (.A(_0457_),
    .B(_0628_),
    .X(_0629_));
 sky130_fd_sc_hd__or3b_1 _1523_ (.A(_0457_),
    .B(_0628_),
    .C_N(_0461_),
    .X(_0630_));
 sky130_fd_sc_hd__nand3_1 _1524_ (.A(_0455_),
    .B(_0459_),
    .C(_0630_),
    .Y(_0631_));
 sky130_fd_sc_hd__a31o_1 _1525_ (.A1(_0455_),
    .A2(_0459_),
    .A3(_0630_),
    .B1(_0453_),
    .X(_0632_));
 sky130_fd_sc_hd__and3_1 _1526_ (.A(_0451_),
    .B(_0454_),
    .C(_0632_),
    .X(_0633_));
 sky130_fd_sc_hd__a21oi_1 _1527_ (.A1(_0451_),
    .A2(_0632_),
    .B1(_0454_),
    .Y(_0634_));
 sky130_fd_sc_hd__or3_1 _1528_ (.A(net183),
    .B(_0633_),
    .C(_0634_),
    .X(_0635_));
 sky130_fd_sc_hd__a22o_1 _1529_ (.A1(\temp_product[39] ),
    .A2(net152),
    .B1(_0625_),
    .B2(_0635_),
    .X(_0278_));
 sky130_fd_sc_hd__xnor2_1 _1530_ (.A(_0453_),
    .B(_0631_),
    .Y(_0636_));
 sky130_fd_sc_hd__or2_1 _1531_ (.A(net183),
    .B(_0636_),
    .X(_0637_));
 sky130_fd_sc_hd__a21o_1 _1532_ (.A1(\temp_product[38] ),
    .A2(net136),
    .B1(net148),
    .X(_0638_));
 sky130_fd_sc_hd__a22o_1 _1533_ (.A1(\temp_product[38] ),
    .A2(net152),
    .B1(_0637_),
    .B2(_0638_),
    .X(_0277_));
 sky130_fd_sc_hd__a21o_1 _1534_ (.A1(\temp_product[37] ),
    .A2(net136),
    .B1(net148),
    .X(_0639_));
 sky130_fd_sc_hd__and3_1 _1535_ (.A(_0455_),
    .B(_0461_),
    .C(_0629_),
    .X(_0640_));
 sky130_fd_sc_hd__a21oi_1 _1536_ (.A1(_0455_),
    .A2(_0629_),
    .B1(_0461_),
    .Y(_0641_));
 sky130_fd_sc_hd__or3_1 _1537_ (.A(net183),
    .B(_0640_),
    .C(_0641_),
    .X(_0642_));
 sky130_fd_sc_hd__a22o_1 _1538_ (.A1(\temp_product[37] ),
    .A2(net152),
    .B1(_0639_),
    .B2(_0642_),
    .X(_0276_));
 sky130_fd_sc_hd__nand2_1 _1539_ (.A(_0457_),
    .B(_0628_),
    .Y(_0643_));
 sky130_fd_sc_hd__a21o_1 _1540_ (.A1(_0629_),
    .A2(_0643_),
    .B1(net183),
    .X(_0644_));
 sky130_fd_sc_hd__a21o_1 _1541_ (.A1(\temp_product[36] ),
    .A2(net136),
    .B1(net148),
    .X(_0645_));
 sky130_fd_sc_hd__a22o_1 _1542_ (.A1(\temp_product[36] ),
    .A2(net152),
    .B1(_0644_),
    .B2(_0645_),
    .X(_0275_));
 sky130_fd_sc_hd__a21o_1 _1543_ (.A1(\temp_product[35] ),
    .A2(net138),
    .B1(net149),
    .X(_0646_));
 sky130_fd_sc_hd__a31o_1 _1544_ (.A1(_0441_),
    .A2(_0445_),
    .A3(_0449_),
    .B1(_0486_),
    .X(_0647_));
 sky130_fd_sc_hd__a21bo_1 _1545_ (.A1(_0447_),
    .A2(_0647_),
    .B1_N(_0446_),
    .X(_0648_));
 sky130_fd_sc_hd__xnor2_1 _1546_ (.A(_0442_),
    .B(_0648_),
    .Y(_0649_));
 sky130_fd_sc_hd__nand2_1 _1547_ (.A(net182),
    .B(_0649_),
    .Y(_0650_));
 sky130_fd_sc_hd__a22o_1 _1548_ (.A1(\temp_product[35] ),
    .A2(net154),
    .B1(_0646_),
    .B2(_0650_),
    .X(_0274_));
 sky130_fd_sc_hd__xnor2_1 _1549_ (.A(_0448_),
    .B(_0647_),
    .Y(_0651_));
 sky130_fd_sc_hd__or2_1 _1550_ (.A(net185),
    .B(_0651_),
    .X(_0652_));
 sky130_fd_sc_hd__a21o_1 _1551_ (.A1(\temp_product[34] ),
    .A2(net140),
    .B1(net150),
    .X(_0653_));
 sky130_fd_sc_hd__a22o_1 _1552_ (.A1(\temp_product[34] ),
    .A2(net155),
    .B1(_0652_),
    .B2(_0653_),
    .X(_0273_));
 sky130_fd_sc_hd__a21o_1 _1553_ (.A1(\temp_product[33] ),
    .A2(net140),
    .B1(net148),
    .X(_0654_));
 sky130_fd_sc_hd__and3_1 _1554_ (.A(_0443_),
    .B(_0449_),
    .C(_0626_),
    .X(_0655_));
 sky130_fd_sc_hd__a21oi_1 _1555_ (.A1(_0443_),
    .A2(_0626_),
    .B1(_0449_),
    .Y(_0656_));
 sky130_fd_sc_hd__or3_1 _1556_ (.A(net183),
    .B(_0655_),
    .C(_0656_),
    .X(_0657_));
 sky130_fd_sc_hd__a22o_1 _1557_ (.A1(\temp_product[33] ),
    .A2(net152),
    .B1(_0654_),
    .B2(_0657_),
    .X(_0272_));
 sky130_fd_sc_hd__or2_1 _1558_ (.A(_0441_),
    .B(_0445_),
    .X(_0658_));
 sky130_fd_sc_hd__a21o_1 _1559_ (.A1(_0626_),
    .A2(_0658_),
    .B1(net183),
    .X(_0659_));
 sky130_fd_sc_hd__a21o_1 _1560_ (.A1(\temp_product[32] ),
    .A2(net137),
    .B1(net148),
    .X(_0660_));
 sky130_fd_sc_hd__a22o_1 _1561_ (.A1(\temp_product[32] ),
    .A2(net152),
    .B1(_0659_),
    .B2(_0660_),
    .X(_0271_));
 sky130_fd_sc_hd__a22o_1 _1562_ (.A1(net127),
    .A2(net169),
    .B1(net138),
    .B2(\temp_product[63] ),
    .X(_0270_));
 sky130_fd_sc_hd__a22o_1 _1563_ (.A1(net126),
    .A2(net169),
    .B1(net139),
    .B2(\temp_product[62] ),
    .X(_0269_));
 sky130_fd_sc_hd__a22o_1 _1564_ (.A1(net125),
    .A2(net169),
    .B1(net139),
    .B2(\temp_product[61] ),
    .X(_0268_));
 sky130_fd_sc_hd__a22o_1 _1565_ (.A1(net124),
    .A2(net170),
    .B1(net142),
    .B2(\temp_product[60] ),
    .X(_0267_));
 sky130_fd_sc_hd__a22o_1 _1566_ (.A1(net122),
    .A2(net170),
    .B1(net143),
    .B2(\temp_product[59] ),
    .X(_0266_));
 sky130_fd_sc_hd__a22o_1 _1567_ (.A1(net121),
    .A2(net170),
    .B1(net143),
    .B2(\temp_product[58] ),
    .X(_0265_));
 sky130_fd_sc_hd__a22o_1 _1568_ (.A1(net120),
    .A2(net170),
    .B1(net142),
    .B2(\temp_product[57] ),
    .X(_0264_));
 sky130_fd_sc_hd__a22o_1 _1569_ (.A1(net119),
    .A2(net170),
    .B1(net142),
    .B2(\temp_product[56] ),
    .X(_0263_));
 sky130_fd_sc_hd__a22o_1 _1570_ (.A1(net118),
    .A2(net170),
    .B1(net141),
    .B2(\temp_product[55] ),
    .X(_0262_));
 sky130_fd_sc_hd__a22o_1 _1571_ (.A1(net117),
    .A2(net171),
    .B1(net141),
    .B2(\temp_product[54] ),
    .X(_0261_));
 sky130_fd_sc_hd__a22o_1 _1572_ (.A1(net116),
    .A2(net170),
    .B1(net142),
    .B2(\temp_product[53] ),
    .X(_0260_));
 sky130_fd_sc_hd__a22o_1 _1573_ (.A1(net115),
    .A2(net171),
    .B1(net141),
    .B2(\temp_product[52] ),
    .X(_0259_));
 sky130_fd_sc_hd__a22o_1 _1574_ (.A1(net114),
    .A2(net171),
    .B1(net143),
    .B2(\temp_product[51] ),
    .X(_0258_));
 sky130_fd_sc_hd__a22o_1 _1575_ (.A1(net113),
    .A2(net171),
    .B1(net141),
    .B2(\temp_product[50] ),
    .X(_0257_));
 sky130_fd_sc_hd__a22o_1 _1576_ (.A1(net111),
    .A2(net171),
    .B1(net141),
    .B2(\temp_product[49] ),
    .X(_0256_));
 sky130_fd_sc_hd__a22o_1 _1577_ (.A1(net110),
    .A2(net171),
    .B1(net141),
    .B2(\temp_product[48] ),
    .X(_0255_));
 sky130_fd_sc_hd__a22o_1 _1578_ (.A1(net109),
    .A2(net169),
    .B1(net138),
    .B2(\temp_product[47] ),
    .X(_0254_));
 sky130_fd_sc_hd__a21o_1 _1579_ (.A1(net108),
    .A2(net169),
    .B1(_0600_),
    .X(_0253_));
 sky130_fd_sc_hd__a22o_1 _1580_ (.A1(net107),
    .A2(net169),
    .B1(net138),
    .B2(\temp_product[45] ),
    .X(_0252_));
 sky130_fd_sc_hd__a22o_1 _1581_ (.A1(net106),
    .A2(net172),
    .B1(net137),
    .B2(\temp_product[44] ),
    .X(_0251_));
 sky130_fd_sc_hd__a22o_1 _1582_ (.A1(net105),
    .A2(net168),
    .B1(net136),
    .B2(\temp_product[43] ),
    .X(_0250_));
 sky130_fd_sc_hd__a22o_1 _1583_ (.A1(net104),
    .A2(net172),
    .B1(net137),
    .B2(\temp_product[42] ),
    .X(_0249_));
 sky130_fd_sc_hd__a22o_1 _1584_ (.A1(net103),
    .A2(net168),
    .B1(net136),
    .B2(\temp_product[41] ),
    .X(_0248_));
 sky130_fd_sc_hd__a22o_1 _1585_ (.A1(net102),
    .A2(net172),
    .B1(net137),
    .B2(\temp_product[40] ),
    .X(_0247_));
 sky130_fd_sc_hd__a22o_1 _1586_ (.A1(net100),
    .A2(net168),
    .B1(net137),
    .B2(\temp_product[39] ),
    .X(_0246_));
 sky130_fd_sc_hd__a22o_1 _1587_ (.A1(net99),
    .A2(net168),
    .B1(net136),
    .B2(\temp_product[38] ),
    .X(_0245_));
 sky130_fd_sc_hd__a22o_1 _1588_ (.A1(net98),
    .A2(net168),
    .B1(net136),
    .B2(\temp_product[37] ),
    .X(_0244_));
 sky130_fd_sc_hd__a22o_1 _1589_ (.A1(net97),
    .A2(net172),
    .B1(net136),
    .B2(\temp_product[36] ),
    .X(_0243_));
 sky130_fd_sc_hd__a22o_1 _1590_ (.A1(net96),
    .A2(net169),
    .B1(net138),
    .B2(\temp_product[35] ),
    .X(_0242_));
 sky130_fd_sc_hd__a22o_1 _1591_ (.A1(net95),
    .A2(net169),
    .B1(net139),
    .B2(\temp_product[34] ),
    .X(_0241_));
 sky130_fd_sc_hd__a22o_1 _1592_ (.A1(net94),
    .A2(net169),
    .B1(net138),
    .B2(\temp_product[33] ),
    .X(_0240_));
 sky130_fd_sc_hd__a22o_1 _1593_ (.A1(net93),
    .A2(net169),
    .B1(net138),
    .B2(\temp_product[32] ),
    .X(_0239_));
 sky130_fd_sc_hd__mux2_1 _1594_ (.A0(\temp_product[31] ),
    .A1(net92),
    .S(net171),
    .X(_0238_));
 sky130_fd_sc_hd__mux2_1 _1595_ (.A0(\temp_product[30] ),
    .A1(net91),
    .S(net168),
    .X(_0237_));
 sky130_fd_sc_hd__mux2_1 _1596_ (.A0(\temp_product[29] ),
    .A1(net89),
    .S(net165),
    .X(_0236_));
 sky130_fd_sc_hd__mux2_1 _1597_ (.A0(\temp_product[28] ),
    .A1(net88),
    .S(net165),
    .X(_0235_));
 sky130_fd_sc_hd__mux2_1 _1598_ (.A0(\temp_product[27] ),
    .A1(net87),
    .S(net166),
    .X(_0234_));
 sky130_fd_sc_hd__mux2_1 _1599_ (.A0(\temp_product[26] ),
    .A1(net86),
    .S(net166),
    .X(_0233_));
 sky130_fd_sc_hd__mux2_1 _1600_ (.A0(\temp_product[25] ),
    .A1(net85),
    .S(net171),
    .X(_0232_));
 sky130_fd_sc_hd__mux2_1 _1601_ (.A0(\temp_product[24] ),
    .A1(net84),
    .S(net171),
    .X(_0231_));
 sky130_fd_sc_hd__mux2_1 _1602_ (.A0(\temp_product[23] ),
    .A1(net83),
    .S(net171),
    .X(_0230_));
 sky130_fd_sc_hd__mux2_1 _1603_ (.A0(\temp_product[22] ),
    .A1(net82),
    .S(net167),
    .X(_0229_));
 sky130_fd_sc_hd__mux2_1 _1604_ (.A0(\temp_product[21] ),
    .A1(net81),
    .S(net167),
    .X(_0228_));
 sky130_fd_sc_hd__mux2_1 _1605_ (.A0(\temp_product[20] ),
    .A1(net80),
    .S(net167),
    .X(_0227_));
 sky130_fd_sc_hd__mux2_1 _1606_ (.A0(\temp_product[19] ),
    .A1(net78),
    .S(net167),
    .X(_0226_));
 sky130_fd_sc_hd__mux2_1 _1607_ (.A0(\temp_product[18] ),
    .A1(net77),
    .S(net166),
    .X(_0225_));
 sky130_fd_sc_hd__mux2_1 _1608_ (.A0(\temp_product[17] ),
    .A1(net76),
    .S(net166),
    .X(_0224_));
 sky130_fd_sc_hd__mux2_1 _1609_ (.A0(\temp_product[16] ),
    .A1(net75),
    .S(net166),
    .X(_0223_));
 sky130_fd_sc_hd__mux2_1 _1610_ (.A0(\temp_product[15] ),
    .A1(net74),
    .S(net166),
    .X(_0222_));
 sky130_fd_sc_hd__mux2_1 _1611_ (.A0(\temp_product[14] ),
    .A1(net73),
    .S(net166),
    .X(_0221_));
 sky130_fd_sc_hd__mux2_1 _1612_ (.A0(\temp_product[13] ),
    .A1(net72),
    .S(net166),
    .X(_0220_));
 sky130_fd_sc_hd__mux2_1 _1613_ (.A0(\temp_product[12] ),
    .A1(net71),
    .S(net166),
    .X(_0219_));
 sky130_fd_sc_hd__mux2_1 _1614_ (.A0(\temp_product[11] ),
    .A1(net70),
    .S(net166),
    .X(_0218_));
 sky130_fd_sc_hd__mux2_1 _1615_ (.A0(\temp_product[10] ),
    .A1(net69),
    .S(net165),
    .X(_0217_));
 sky130_fd_sc_hd__mux2_1 _1616_ (.A0(\temp_product[9] ),
    .A1(net131),
    .S(net165),
    .X(_0216_));
 sky130_fd_sc_hd__mux2_1 _1617_ (.A0(\temp_product[8] ),
    .A1(net130),
    .S(net165),
    .X(_0215_));
 sky130_fd_sc_hd__mux2_1 _1618_ (.A0(\temp_product[7] ),
    .A1(net129),
    .S(net165),
    .X(_0214_));
 sky130_fd_sc_hd__mux2_1 _1619_ (.A0(\temp_product[6] ),
    .A1(net128),
    .S(net165),
    .X(_0213_));
 sky130_fd_sc_hd__mux2_1 _1620_ (.A0(\temp_product[5] ),
    .A1(net123),
    .S(net165),
    .X(_0212_));
 sky130_fd_sc_hd__mux2_1 _1621_ (.A0(\temp_product[4] ),
    .A1(net112),
    .S(net165),
    .X(_0211_));
 sky130_fd_sc_hd__mux2_1 _1622_ (.A0(\temp_product[3] ),
    .A1(net101),
    .S(net165),
    .X(_0210_));
 sky130_fd_sc_hd__mux2_1 _1623_ (.A0(\temp_product[2] ),
    .A1(net90),
    .S(net167),
    .X(_0209_));
 sky130_fd_sc_hd__mux2_1 _1624_ (.A0(\temp_product[1] ),
    .A1(net79),
    .S(net167),
    .X(_0208_));
 sky130_fd_sc_hd__mux2_1 _1625_ (.A0(\temp_product[0] ),
    .A1(net68),
    .S(net168),
    .X(_0207_));
 sky130_fd_sc_hd__a21o_1 _1626_ (.A1(\count[5] ),
    .A2(_0668_),
    .B1(net203),
    .X(_0206_));
 sky130_fd_sc_hd__nand2_1 _1627_ (.A(\count[4] ),
    .B(_0667_),
    .Y(_0661_));
 sky130_fd_sc_hd__a21oi_1 _1628_ (.A1(_0668_),
    .A2(_0661_),
    .B1(_0674_),
    .Y(_0205_));
 sky130_fd_sc_hd__nand2_1 _1629_ (.A(\count[3] ),
    .B(_0666_),
    .Y(_0662_));
 sky130_fd_sc_hd__a21oi_1 _1630_ (.A1(_0667_),
    .A2(_0662_),
    .B1(_0674_),
    .Y(_0204_));
 sky130_fd_sc_hd__nand2_1 _1631_ (.A(\count[2] ),
    .B(_0665_),
    .Y(_0663_));
 sky130_fd_sc_hd__a21oi_1 _1632_ (.A1(_0666_),
    .A2(_0663_),
    .B1(_0674_),
    .Y(_0203_));
 sky130_fd_sc_hd__nand2_1 _1633_ (.A(\count[1] ),
    .B(\count[0] ),
    .Y(_0664_));
 sky130_fd_sc_hd__a21oi_1 _1634_ (.A1(_0665_),
    .A2(_0664_),
    .B1(_0674_),
    .Y(_0202_));
 sky130_fd_sc_hd__nor2_1 _1635_ (.A(\count[0] ),
    .B(_0674_),
    .Y(_0201_));
 sky130_fd_sc_hd__mux2_1 _1636_ (.A0(\b[31] ),
    .A1(net57),
    .S(net202),
    .X(_0200_));
 sky130_fd_sc_hd__o21ba_1 _1637_ (.A1(net67),
    .A2(net184),
    .B1_N(net204),
    .X(_0199_));
 sky130_fd_sc_hd__inv_2 _1638_ (.A(net221),
    .Y(_0001_));
 sky130_fd_sc_hd__inv_2 _1639_ (.A(net223),
    .Y(_0002_));
 sky130_fd_sc_hd__inv_2 _1640_ (.A(net223),
    .Y(_0003_));
 sky130_fd_sc_hd__inv_2 _1641_ (.A(net221),
    .Y(_0004_));
 sky130_fd_sc_hd__inv_2 _1642_ (.A(net221),
    .Y(_0005_));
 sky130_fd_sc_hd__inv_2 _1643_ (.A(net223),
    .Y(_0006_));
 sky130_fd_sc_hd__inv_2 _1644_ (.A(net223),
    .Y(_0007_));
 sky130_fd_sc_hd__inv_2 _1645_ (.A(net224),
    .Y(_0008_));
 sky130_fd_sc_hd__inv_2 _1646_ (.A(net210),
    .Y(_0009_));
 sky130_fd_sc_hd__inv_2 _1647_ (.A(net210),
    .Y(_0010_));
 sky130_fd_sc_hd__inv_2 _1648_ (.A(net206),
    .Y(_0011_));
 sky130_fd_sc_hd__inv_2 _1649_ (.A(net208),
    .Y(_0012_));
 sky130_fd_sc_hd__inv_2 _1650_ (.A(net208),
    .Y(_0013_));
 sky130_fd_sc_hd__inv_2 _1651_ (.A(net208),
    .Y(_0014_));
 sky130_fd_sc_hd__inv_2 _1652_ (.A(net206),
    .Y(_0015_));
 sky130_fd_sc_hd__inv_2 _1653_ (.A(net208),
    .Y(_0016_));
 sky130_fd_sc_hd__inv_2 _1654_ (.A(net208),
    .Y(_0017_));
 sky130_fd_sc_hd__inv_2 _1655_ (.A(net208),
    .Y(_0018_));
 sky130_fd_sc_hd__inv_2 _1656_ (.A(net214),
    .Y(_0019_));
 sky130_fd_sc_hd__inv_2 _1657_ (.A(net216),
    .Y(_0020_));
 sky130_fd_sc_hd__inv_2 _1658_ (.A(net216),
    .Y(_0021_));
 sky130_fd_sc_hd__inv_2 _1659_ (.A(net216),
    .Y(_0022_));
 sky130_fd_sc_hd__inv_2 _1660_ (.A(net216),
    .Y(_0023_));
 sky130_fd_sc_hd__inv_2 _1661_ (.A(net214),
    .Y(_0024_));
 sky130_fd_sc_hd__inv_2 _1662_ (.A(net216),
    .Y(_0025_));
 sky130_fd_sc_hd__inv_2 _1663_ (.A(net218),
    .Y(_0026_));
 sky130_fd_sc_hd__inv_2 _1664_ (.A(net218),
    .Y(_0027_));
 sky130_fd_sc_hd__inv_2 _1665_ (.A(net218),
    .Y(_0028_));
 sky130_fd_sc_hd__inv_2 _1666_ (.A(net218),
    .Y(_0029_));
 sky130_fd_sc_hd__inv_2 _1667_ (.A(net218),
    .Y(_0030_));
 sky130_fd_sc_hd__inv_2 _1668_ (.A(net227),
    .Y(_0031_));
 sky130_fd_sc_hd__inv_2 _1669_ (.A(net227),
    .Y(_0032_));
 sky130_fd_sc_hd__inv_2 _1670_ (.A(net227),
    .Y(_0033_));
 sky130_fd_sc_hd__inv_2 _1671_ (.A(net214),
    .Y(_0034_));
 sky130_fd_sc_hd__inv_2 _1672_ (.A(net214),
    .Y(_0035_));
 sky130_fd_sc_hd__inv_2 _1673_ (.A(net208),
    .Y(_0036_));
 sky130_fd_sc_hd__inv_2 _1674_ (.A(net210),
    .Y(_0037_));
 sky130_fd_sc_hd__inv_2 _1675_ (.A(net224),
    .Y(_0038_));
 sky130_fd_sc_hd__inv_2 _1676_ (.A(net227),
    .Y(_0039_));
 sky130_fd_sc_hd__inv_2 _1677_ (.A(net230),
    .Y(_0040_));
 sky130_fd_sc_hd__inv_2 _1678_ (.A(net230),
    .Y(_0041_));
 sky130_fd_sc_hd__inv_2 _1679_ (.A(net230),
    .Y(_0042_));
 sky130_fd_sc_hd__inv_2 _1680_ (.A(net230),
    .Y(_0043_));
 sky130_fd_sc_hd__inv_2 _1681_ (.A(net224),
    .Y(_0044_));
 sky130_fd_sc_hd__inv_2 _1682_ (.A(net221),
    .Y(_0045_));
 sky130_fd_sc_hd__inv_2 _1683_ (.A(net224),
    .Y(_0046_));
 sky130_fd_sc_hd__inv_2 _1684_ (.A(net225),
    .Y(_0047_));
 sky130_fd_sc_hd__inv_2 _1685_ (.A(net225),
    .Y(_0048_));
 sky130_fd_sc_hd__inv_2 _1686_ (.A(net224),
    .Y(_0049_));
 sky130_fd_sc_hd__inv_2 _1687_ (.A(net225),
    .Y(_0050_));
 sky130_fd_sc_hd__inv_2 _1688_ (.A(net225),
    .Y(_0051_));
 sky130_fd_sc_hd__inv_2 _1689_ (.A(net225),
    .Y(_0052_));
 sky130_fd_sc_hd__inv_2 _1690_ (.A(net225),
    .Y(_0053_));
 sky130_fd_sc_hd__inv_2 _1691_ (.A(net230),
    .Y(_0054_));
 sky130_fd_sc_hd__inv_2 _1692_ (.A(net230),
    .Y(_0055_));
 sky130_fd_sc_hd__inv_2 _1693_ (.A(net227),
    .Y(_0056_));
 sky130_fd_sc_hd__inv_2 _1694_ (.A(net227),
    .Y(_0057_));
 sky130_fd_sc_hd__inv_2 _1695_ (.A(net227),
    .Y(_0058_));
 sky130_fd_sc_hd__inv_2 _1696_ (.A(net228),
    .Y(_0059_));
 sky130_fd_sc_hd__inv_2 _1697_ (.A(net228),
    .Y(_0060_));
 sky130_fd_sc_hd__inv_2 _1698_ (.A(net232),
    .Y(_0061_));
 sky130_fd_sc_hd__inv_2 _1699_ (.A(net228),
    .Y(_0062_));
 sky130_fd_sc_hd__inv_2 _1700_ (.A(net232),
    .Y(_0063_));
 sky130_fd_sc_hd__inv_2 _1701_ (.A(net232),
    .Y(_0064_));
 sky130_fd_sc_hd__inv_2 _1702_ (.A(net232),
    .Y(_0065_));
 sky130_fd_sc_hd__inv_2 _1703_ (.A(net232),
    .Y(_0066_));
 sky130_fd_sc_hd__inv_2 _1704_ (.A(net232),
    .Y(_0067_));
 sky130_fd_sc_hd__inv_2 _1705_ (.A(net233),
    .Y(_0068_));
 sky130_fd_sc_hd__inv_2 _1706_ (.A(net230),
    .Y(_0069_));
 sky130_fd_sc_hd__inv_2 _1707_ (.A(net230),
    .Y(_0070_));
 sky130_fd_sc_hd__inv_2 _1708_ (.A(net230),
    .Y(_0071_));
 sky130_fd_sc_hd__inv_2 _1709_ (.A(net223),
    .Y(_0072_));
 sky130_fd_sc_hd__inv_2 _1710_ (.A(net229),
    .Y(_0073_));
 sky130_fd_sc_hd__inv_2 _1711_ (.A(net229),
    .Y(_0074_));
 sky130_fd_sc_hd__inv_2 _1712_ (.A(net231),
    .Y(_0075_));
 sky130_fd_sc_hd__inv_2 _1713_ (.A(net224),
    .Y(_0076_));
 sky130_fd_sc_hd__inv_2 _1714_ (.A(net222),
    .Y(_0077_));
 sky130_fd_sc_hd__inv_2 _1715_ (.A(net222),
    .Y(_0078_));
 sky130_fd_sc_hd__inv_2 _1716_ (.A(net223),
    .Y(_0079_));
 sky130_fd_sc_hd__inv_2 _1717_ (.A(net225),
    .Y(_0080_));
 sky130_fd_sc_hd__inv_2 _1718_ (.A(net224),
    .Y(_0081_));
 sky130_fd_sc_hd__inv_2 _1719_ (.A(net226),
    .Y(_0082_));
 sky130_fd_sc_hd__inv_2 _1720_ (.A(net225),
    .Y(_0083_));
 sky130_fd_sc_hd__inv_2 _1721_ (.A(net226),
    .Y(_0084_));
 sky130_fd_sc_hd__inv_2 _1722_ (.A(net230),
    .Y(_0085_));
 sky130_fd_sc_hd__inv_2 _1723_ (.A(net226),
    .Y(_0086_));
 sky130_fd_sc_hd__inv_2 _1724_ (.A(net231),
    .Y(_0087_));
 sky130_fd_sc_hd__inv_2 _1725_ (.A(net229),
    .Y(_0088_));
 sky130_fd_sc_hd__inv_2 _1726_ (.A(net227),
    .Y(_0089_));
 sky130_fd_sc_hd__inv_2 _1727_ (.A(net227),
    .Y(_0090_));
 sky130_fd_sc_hd__inv_2 _1728_ (.A(net228),
    .Y(_0091_));
 sky130_fd_sc_hd__inv_2 _1729_ (.A(net229),
    .Y(_0092_));
 sky130_fd_sc_hd__inv_2 _1730_ (.A(net232),
    .Y(_0093_));
 sky130_fd_sc_hd__inv_2 _1731_ (.A(net228),
    .Y(_0094_));
 sky130_fd_sc_hd__inv_2 _1732_ (.A(net232),
    .Y(_0095_));
 sky130_fd_sc_hd__inv_2 _1733_ (.A(net232),
    .Y(_0096_));
 sky130_fd_sc_hd__inv_2 _1734_ (.A(net232),
    .Y(_0097_));
 sky130_fd_sc_hd__inv_2 _1735_ (.A(net233),
    .Y(_0098_));
 sky130_fd_sc_hd__inv_2 _1736_ (.A(net233),
    .Y(_0099_));
 sky130_fd_sc_hd__inv_2 _1737_ (.A(net233),
    .Y(_0100_));
 sky130_fd_sc_hd__inv_2 _1738_ (.A(net231),
    .Y(_0101_));
 sky130_fd_sc_hd__inv_2 _1739_ (.A(net231),
    .Y(_0102_));
 sky130_fd_sc_hd__inv_2 _1740_ (.A(net231),
    .Y(_0103_));
 sky130_fd_sc_hd__inv_2 _1741_ (.A(net210),
    .Y(_0104_));
 sky130_fd_sc_hd__inv_2 _1742_ (.A(net211),
    .Y(_0105_));
 sky130_fd_sc_hd__inv_2 _1743_ (.A(net210),
    .Y(_0106_));
 sky130_fd_sc_hd__inv_2 _1744_ (.A(net207),
    .Y(_0107_));
 sky130_fd_sc_hd__inv_2 _1745_ (.A(net207),
    .Y(_0108_));
 sky130_fd_sc_hd__inv_2 _1746_ (.A(net206),
    .Y(_0109_));
 sky130_fd_sc_hd__inv_2 _1747_ (.A(net206),
    .Y(_0110_));
 sky130_fd_sc_hd__inv_2 _1748_ (.A(net208),
    .Y(_0111_));
 sky130_fd_sc_hd__inv_2 _1749_ (.A(net208),
    .Y(_0112_));
 sky130_fd_sc_hd__inv_2 _1750_ (.A(net214),
    .Y(_0113_));
 sky130_fd_sc_hd__inv_2 _1751_ (.A(net214),
    .Y(_0114_));
 sky130_fd_sc_hd__inv_2 _1752_ (.A(net214),
    .Y(_0115_));
 sky130_fd_sc_hd__inv_2 _1753_ (.A(net214),
    .Y(_0116_));
 sky130_fd_sc_hd__inv_2 _1754_ (.A(net214),
    .Y(_0117_));
 sky130_fd_sc_hd__inv_2 _1755_ (.A(net216),
    .Y(_0118_));
 sky130_fd_sc_hd__inv_2 _1756_ (.A(net216),
    .Y(_0119_));
 sky130_fd_sc_hd__inv_2 _1757_ (.A(net214),
    .Y(_0120_));
 sky130_fd_sc_hd__inv_2 _1758_ (.A(net215),
    .Y(_0121_));
 sky130_fd_sc_hd__inv_2 _1759_ (.A(net216),
    .Y(_0122_));
 sky130_fd_sc_hd__inv_2 _1760_ (.A(net217),
    .Y(_0123_));
 sky130_fd_sc_hd__inv_2 _1761_ (.A(net218),
    .Y(_0124_));
 sky130_fd_sc_hd__inv_2 _1762_ (.A(net218),
    .Y(_0125_));
 sky130_fd_sc_hd__inv_2 _1763_ (.A(net220),
    .Y(_0126_));
 sky130_fd_sc_hd__inv_2 _1764_ (.A(net219),
    .Y(_0127_));
 sky130_fd_sc_hd__inv_2 _1765_ (.A(net219),
    .Y(_0128_));
 sky130_fd_sc_hd__inv_2 _1766_ (.A(net219),
    .Y(_0129_));
 sky130_fd_sc_hd__inv_2 _1767_ (.A(net219),
    .Y(_0130_));
 sky130_fd_sc_hd__inv_2 _1768_ (.A(net209),
    .Y(_0131_));
 sky130_fd_sc_hd__inv_2 _1769_ (.A(net212),
    .Y(_0132_));
 sky130_fd_sc_hd__inv_2 _1770_ (.A(net212),
    .Y(_0133_));
 sky130_fd_sc_hd__inv_2 _1771_ (.A(net212),
    .Y(_0134_));
 sky130_fd_sc_hd__inv_2 _1772_ (.A(net212),
    .Y(_0135_));
 sky130_fd_sc_hd__inv_2 _1773_ (.A(net221),
    .Y(_0136_));
 sky130_fd_sc_hd__inv_2 _1774_ (.A(net222),
    .Y(_0137_));
 sky130_fd_sc_hd__inv_2 _1775_ (.A(net224),
    .Y(_0138_));
 sky130_fd_sc_hd__inv_2 _1776_ (.A(net224),
    .Y(_0139_));
 sky130_fd_sc_hd__inv_2 _1777_ (.A(net211),
    .Y(_0140_));
 sky130_fd_sc_hd__inv_2 _1778_ (.A(net210),
    .Y(_0141_));
 sky130_fd_sc_hd__inv_2 _1779_ (.A(net210),
    .Y(_0142_));
 sky130_fd_sc_hd__inv_2 _1780_ (.A(net207),
    .Y(_0143_));
 sky130_fd_sc_hd__inv_2 _1781_ (.A(net207),
    .Y(_0144_));
 sky130_fd_sc_hd__inv_2 _1782_ (.A(net207),
    .Y(_0145_));
 sky130_fd_sc_hd__inv_2 _1783_ (.A(net206),
    .Y(_0146_));
 sky130_fd_sc_hd__inv_2 _1784_ (.A(net206),
    .Y(_0147_));
 sky130_fd_sc_hd__inv_2 _1785_ (.A(net206),
    .Y(_0148_));
 sky130_fd_sc_hd__inv_2 _1786_ (.A(net206),
    .Y(_0149_));
 sky130_fd_sc_hd__inv_2 _1787_ (.A(net206),
    .Y(_0150_));
 sky130_fd_sc_hd__inv_2 _1788_ (.A(net207),
    .Y(_0151_));
 sky130_fd_sc_hd__inv_2 _1789_ (.A(net210),
    .Y(_0152_));
 sky130_fd_sc_hd__inv_2 _1790_ (.A(net210),
    .Y(_0153_));
 sky130_fd_sc_hd__inv_2 _1791_ (.A(net211),
    .Y(_0154_));
 sky130_fd_sc_hd__inv_2 _1792_ (.A(net211),
    .Y(_0155_));
 sky130_fd_sc_hd__inv_2 _1793_ (.A(net211),
    .Y(_0156_));
 sky130_fd_sc_hd__inv_2 _1794_ (.A(net221),
    .Y(_0157_));
 sky130_fd_sc_hd__inv_2 _1795_ (.A(net221),
    .Y(_0158_));
 sky130_fd_sc_hd__inv_2 _1796_ (.A(net224),
    .Y(_0159_));
 sky130_fd_sc_hd__inv_2 _1797_ (.A(net222),
    .Y(_0160_));
 sky130_fd_sc_hd__inv_2 _1798_ (.A(net222),
    .Y(_0161_));
 sky130_fd_sc_hd__inv_2 _1799_ (.A(net222),
    .Y(_0162_));
 sky130_fd_sc_hd__inv_2 _1800_ (.A(net222),
    .Y(_0163_));
 sky130_fd_sc_hd__inv_2 _1801_ (.A(net221),
    .Y(_0164_));
 sky130_fd_sc_hd__inv_2 _1802_ (.A(net221),
    .Y(_0165_));
 sky130_fd_sc_hd__inv_2 _1803_ (.A(net221),
    .Y(_0166_));
 sky130_fd_sc_hd__inv_2 _1804_ (.A(net211),
    .Y(_0167_));
 sky130_fd_sc_hd__inv_2 _1805_ (.A(net211),
    .Y(_0168_));
 sky130_fd_sc_hd__inv_2 _1806_ (.A(net210),
    .Y(_0169_));
 sky130_fd_sc_hd__inv_2 _1807_ (.A(net207),
    .Y(_0170_));
 sky130_fd_sc_hd__inv_2 _1808_ (.A(net209),
    .Y(_0171_));
 sky130_fd_sc_hd__inv_2 _1809_ (.A(net206),
    .Y(_0172_));
 sky130_fd_sc_hd__inv_2 _1810_ (.A(net209),
    .Y(_0173_));
 sky130_fd_sc_hd__inv_2 _1811_ (.A(net208),
    .Y(_0174_));
 sky130_fd_sc_hd__inv_2 _1812_ (.A(net209),
    .Y(_0175_));
 sky130_fd_sc_hd__inv_2 _1813_ (.A(net209),
    .Y(_0176_));
 sky130_fd_sc_hd__inv_2 _1814_ (.A(net215),
    .Y(_0177_));
 sky130_fd_sc_hd__inv_2 _1815_ (.A(net215),
    .Y(_0178_));
 sky130_fd_sc_hd__inv_2 _1816_ (.A(net217),
    .Y(_0179_));
 sky130_fd_sc_hd__inv_2 _1817_ (.A(net216),
    .Y(_0180_));
 sky130_fd_sc_hd__inv_2 _1818_ (.A(net216),
    .Y(_0181_));
 sky130_fd_sc_hd__inv_2 _1819_ (.A(net217),
    .Y(_0182_));
 sky130_fd_sc_hd__inv_2 _1820_ (.A(net215),
    .Y(_0183_));
 sky130_fd_sc_hd__inv_2 _1821_ (.A(net217),
    .Y(_0184_));
 sky130_fd_sc_hd__inv_2 _1822_ (.A(net217),
    .Y(_0185_));
 sky130_fd_sc_hd__inv_2 _1823_ (.A(net218),
    .Y(_0186_));
 sky130_fd_sc_hd__inv_2 _1824_ (.A(net218),
    .Y(_0187_));
 sky130_fd_sc_hd__inv_2 _1825_ (.A(net218),
    .Y(_0188_));
 sky130_fd_sc_hd__inv_2 _1826_ (.A(net227),
    .Y(_0189_));
 sky130_fd_sc_hd__inv_2 _1827_ (.A(net219),
    .Y(_0190_));
 sky130_fd_sc_hd__inv_2 _1828_ (.A(net219),
    .Y(_0191_));
 sky130_fd_sc_hd__inv_2 _1829_ (.A(net219),
    .Y(_0192_));
 sky130_fd_sc_hd__inv_2 _1830_ (.A(net219),
    .Y(_0193_));
 sky130_fd_sc_hd__inv_2 _1831_ (.A(net215),
    .Y(_0194_));
 sky130_fd_sc_hd__inv_2 _1832_ (.A(net212),
    .Y(_0195_));
 sky130_fd_sc_hd__inv_2 _1833_ (.A(net212),
    .Y(_0196_));
 sky130_fd_sc_hd__inv_2 _1834_ (.A(net212),
    .Y(_0197_));
 sky130_fd_sc_hd__inv_2 _1835_ (.A(net219),
    .Y(_0198_));
 sky130_fd_sc_hd__dfrtp_1 _1836_ (.CLK(clknet_4_7_0_clk),
    .D(_0199_),
    .RESET_B(_0000_),
    .Q(net67));
 sky130_fd_sc_hd__dfrtp_1 _1837_ (.CLK(clknet_4_4_0_clk),
    .D(_0200_),
    .RESET_B(_0001_),
    .Q(\b[31] ));
 sky130_fd_sc_hd__dfrtp_1 _1838_ (.CLK(clknet_4_4_0_clk),
    .D(_0201_),
    .RESET_B(_0002_),
    .Q(\count[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1839_ (.CLK(clknet_4_6_0_clk),
    .D(_0202_),
    .RESET_B(_0003_),
    .Q(\count[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1840_ (.CLK(clknet_4_4_0_clk),
    .D(_0203_),
    .RESET_B(_0004_),
    .Q(\count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1841_ (.CLK(clknet_4_4_0_clk),
    .D(_0204_),
    .RESET_B(_0005_),
    .Q(\count[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1842_ (.CLK(clknet_4_6_0_clk),
    .D(_0205_),
    .RESET_B(_0006_),
    .Q(\count[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1843_ (.CLK(clknet_4_6_0_clk),
    .D(_0206_),
    .RESET_B(_0007_),
    .Q(\count[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1844_ (.CLK(clknet_4_5_0_clk),
    .D(_0207_),
    .RESET_B(_0008_),
    .Q(net68));
 sky130_fd_sc_hd__dfrtp_1 _1845_ (.CLK(clknet_4_1_0_clk),
    .D(_0208_),
    .RESET_B(_0009_),
    .Q(net79));
 sky130_fd_sc_hd__dfrtp_1 _1846_ (.CLK(clknet_4_1_0_clk),
    .D(_0209_),
    .RESET_B(_0010_),
    .Q(net90));
 sky130_fd_sc_hd__dfrtp_1 _1847_ (.CLK(clknet_4_0_0_clk),
    .D(_0210_),
    .RESET_B(_0011_),
    .Q(net101));
 sky130_fd_sc_hd__dfrtp_1 _1848_ (.CLK(clknet_4_2_0_clk),
    .D(_0211_),
    .RESET_B(_0012_),
    .Q(net112));
 sky130_fd_sc_hd__dfrtp_1 _1849_ (.CLK(clknet_4_2_0_clk),
    .D(_0212_),
    .RESET_B(_0013_),
    .Q(net123));
 sky130_fd_sc_hd__dfrtp_1 _1850_ (.CLK(clknet_4_2_0_clk),
    .D(_0213_),
    .RESET_B(_0014_),
    .Q(net128));
 sky130_fd_sc_hd__dfrtp_1 _1851_ (.CLK(clknet_4_0_0_clk),
    .D(_0214_),
    .RESET_B(_0015_),
    .Q(net129));
 sky130_fd_sc_hd__dfrtp_1 _1852_ (.CLK(clknet_4_2_0_clk),
    .D(_0215_),
    .RESET_B(_0016_),
    .Q(net130));
 sky130_fd_sc_hd__dfrtp_1 _1853_ (.CLK(clknet_4_2_0_clk),
    .D(_0216_),
    .RESET_B(_0017_),
    .Q(net131));
 sky130_fd_sc_hd__dfrtp_1 _1854_ (.CLK(clknet_4_2_0_clk),
    .D(_0217_),
    .RESET_B(_0018_),
    .Q(net69));
 sky130_fd_sc_hd__dfrtp_1 _1855_ (.CLK(clknet_4_8_0_clk),
    .D(_0218_),
    .RESET_B(_0019_),
    .Q(net70));
 sky130_fd_sc_hd__dfrtp_1 _1856_ (.CLK(clknet_4_8_0_clk),
    .D(_0219_),
    .RESET_B(_0020_),
    .Q(net71));
 sky130_fd_sc_hd__dfrtp_1 _1857_ (.CLK(clknet_4_10_0_clk),
    .D(_0220_),
    .RESET_B(_0021_),
    .Q(net72));
 sky130_fd_sc_hd__dfrtp_1 _1858_ (.CLK(clknet_4_10_0_clk),
    .D(_0221_),
    .RESET_B(_0022_),
    .Q(net73));
 sky130_fd_sc_hd__dfrtp_1 _1859_ (.CLK(clknet_4_10_0_clk),
    .D(_0222_),
    .RESET_B(_0023_),
    .Q(net74));
 sky130_fd_sc_hd__dfrtp_1 _1860_ (.CLK(clknet_4_8_0_clk),
    .D(_0223_),
    .RESET_B(_0024_),
    .Q(net75));
 sky130_fd_sc_hd__dfrtp_1 _1861_ (.CLK(clknet_4_10_0_clk),
    .D(_0224_),
    .RESET_B(_0025_),
    .Q(net76));
 sky130_fd_sc_hd__dfrtp_1 _1862_ (.CLK(clknet_4_10_0_clk),
    .D(_0225_),
    .RESET_B(_0026_),
    .Q(net77));
 sky130_fd_sc_hd__dfrtp_1 _1863_ (.CLK(clknet_4_11_0_clk),
    .D(_0226_),
    .RESET_B(_0027_),
    .Q(net78));
 sky130_fd_sc_hd__dfrtp_1 _1864_ (.CLK(clknet_4_11_0_clk),
    .D(_0227_),
    .RESET_B(_0028_),
    .Q(net80));
 sky130_fd_sc_hd__dfrtp_1 _1865_ (.CLK(clknet_4_11_0_clk),
    .D(_0228_),
    .RESET_B(_0029_),
    .Q(net81));
 sky130_fd_sc_hd__dfrtp_1 _1866_ (.CLK(clknet_4_11_0_clk),
    .D(_0229_),
    .RESET_B(_0030_),
    .Q(net82));
 sky130_fd_sc_hd__dfrtp_1 _1867_ (.CLK(clknet_4_14_0_clk),
    .D(_0230_),
    .RESET_B(_0031_),
    .Q(net83));
 sky130_fd_sc_hd__dfrtp_1 _1868_ (.CLK(clknet_4_14_0_clk),
    .D(_0231_),
    .RESET_B(_0032_),
    .Q(net84));
 sky130_fd_sc_hd__dfrtp_1 _1869_ (.CLK(clknet_4_11_0_clk),
    .D(_0232_),
    .RESET_B(_0033_),
    .Q(net85));
 sky130_fd_sc_hd__dfrtp_1 _1870_ (.CLK(clknet_4_8_0_clk),
    .D(_0233_),
    .RESET_B(_0034_),
    .Q(net86));
 sky130_fd_sc_hd__dfrtp_1 _1871_ (.CLK(clknet_4_2_0_clk),
    .D(_0234_),
    .RESET_B(_0035_),
    .Q(net87));
 sky130_fd_sc_hd__dfrtp_1 _1872_ (.CLK(clknet_4_2_0_clk),
    .D(_0235_),
    .RESET_B(_0036_),
    .Q(net88));
 sky130_fd_sc_hd__dfrtp_1 _1873_ (.CLK(clknet_4_1_0_clk),
    .D(_0236_),
    .RESET_B(_0037_),
    .Q(net89));
 sky130_fd_sc_hd__dfrtp_1 _1874_ (.CLK(clknet_4_5_0_clk),
    .D(_0237_),
    .RESET_B(_0038_),
    .Q(net91));
 sky130_fd_sc_hd__dfrtp_1 _1875_ (.CLK(clknet_4_14_0_clk),
    .D(_0238_),
    .RESET_B(_0039_),
    .Q(net92));
 sky130_fd_sc_hd__dfrtp_1 _1876_ (.CLK(clknet_4_12_0_clk),
    .D(_0239_),
    .RESET_B(_0040_),
    .Q(net93));
 sky130_fd_sc_hd__dfrtp_1 _1877_ (.CLK(clknet_4_12_0_clk),
    .D(_0240_),
    .RESET_B(_0041_),
    .Q(net94));
 sky130_fd_sc_hd__dfrtp_1 _1878_ (.CLK(clknet_4_13_0_clk),
    .D(_0241_),
    .RESET_B(_0042_),
    .Q(net95));
 sky130_fd_sc_hd__dfrtp_1 _1879_ (.CLK(clknet_4_12_0_clk),
    .D(_0242_),
    .RESET_B(_0043_),
    .Q(net96));
 sky130_fd_sc_hd__dfrtp_1 _1880_ (.CLK(clknet_4_5_0_clk),
    .D(_0243_),
    .RESET_B(_0044_),
    .Q(net97));
 sky130_fd_sc_hd__dfrtp_1 _1881_ (.CLK(clknet_4_4_0_clk),
    .D(_0244_),
    .RESET_B(_0045_),
    .Q(net98));
 sky130_fd_sc_hd__dfrtp_1 _1882_ (.CLK(clknet_4_5_0_clk),
    .D(_0245_),
    .RESET_B(_0046_),
    .Q(net99));
 sky130_fd_sc_hd__dfrtp_1 _1883_ (.CLK(clknet_4_7_0_clk),
    .D(_0246_),
    .RESET_B(_0047_),
    .Q(net100));
 sky130_fd_sc_hd__dfrtp_1 _1884_ (.CLK(clknet_4_7_0_clk),
    .D(_0247_),
    .RESET_B(_0048_),
    .Q(net102));
 sky130_fd_sc_hd__dfrtp_1 _1885_ (.CLK(clknet_4_5_0_clk),
    .D(_0248_),
    .RESET_B(_0049_),
    .Q(net103));
 sky130_fd_sc_hd__dfrtp_1 _1886_ (.CLK(clknet_4_7_0_clk),
    .D(_0249_),
    .RESET_B(_0050_),
    .Q(net104));
 sky130_fd_sc_hd__dfrtp_1 _1887_ (.CLK(clknet_4_5_0_clk),
    .D(_0250_),
    .RESET_B(_0051_),
    .Q(net105));
 sky130_fd_sc_hd__dfrtp_1 _1888_ (.CLK(clknet_4_7_0_clk),
    .D(_0251_),
    .RESET_B(_0052_),
    .Q(net106));
 sky130_fd_sc_hd__dfrtp_1 _1889_ (.CLK(clknet_4_7_0_clk),
    .D(_0252_),
    .RESET_B(_0053_),
    .Q(net107));
 sky130_fd_sc_hd__dfrtp_1 _1890_ (.CLK(clknet_4_13_0_clk),
    .D(_0253_),
    .RESET_B(_0054_),
    .Q(net108));
 sky130_fd_sc_hd__dfrtp_1 _1891_ (.CLK(clknet_4_13_0_clk),
    .D(_0254_),
    .RESET_B(_0055_),
    .Q(net109));
 sky130_fd_sc_hd__dfrtp_1 _1892_ (.CLK(clknet_4_14_0_clk),
    .D(_0255_),
    .RESET_B(_0056_),
    .Q(net110));
 sky130_fd_sc_hd__dfrtp_1 _1893_ (.CLK(clknet_4_14_0_clk),
    .D(_0256_),
    .RESET_B(_0057_),
    .Q(net111));
 sky130_fd_sc_hd__dfrtp_1 _1894_ (.CLK(clknet_4_14_0_clk),
    .D(_0257_),
    .RESET_B(_0058_),
    .Q(net113));
 sky130_fd_sc_hd__dfrtp_1 _1895_ (.CLK(clknet_4_14_0_clk),
    .D(_0258_),
    .RESET_B(_0059_),
    .Q(net114));
 sky130_fd_sc_hd__dfrtp_1 _1896_ (.CLK(clknet_4_14_0_clk),
    .D(_0259_),
    .RESET_B(_0060_),
    .Q(net115));
 sky130_fd_sc_hd__dfrtp_1 _1897_ (.CLK(clknet_4_15_0_clk),
    .D(_0260_),
    .RESET_B(_0061_),
    .Q(net116));
 sky130_fd_sc_hd__dfrtp_1 _1898_ (.CLK(clknet_4_15_0_clk),
    .D(_0261_),
    .RESET_B(_0062_),
    .Q(net117));
 sky130_fd_sc_hd__dfrtp_1 _1899_ (.CLK(clknet_4_15_0_clk),
    .D(_0262_),
    .RESET_B(_0063_),
    .Q(net118));
 sky130_fd_sc_hd__dfrtp_1 _1900_ (.CLK(clknet_4_15_0_clk),
    .D(_0263_),
    .RESET_B(_0064_),
    .Q(net119));
 sky130_fd_sc_hd__dfrtp_1 _1901_ (.CLK(clknet_4_15_0_clk),
    .D(_0264_),
    .RESET_B(_0065_),
    .Q(net120));
 sky130_fd_sc_hd__dfrtp_1 _1902_ (.CLK(clknet_4_15_0_clk),
    .D(_0265_),
    .RESET_B(_0066_),
    .Q(net121));
 sky130_fd_sc_hd__dfrtp_1 _1903_ (.CLK(clknet_4_15_0_clk),
    .D(_0266_),
    .RESET_B(_0067_),
    .Q(net122));
 sky130_fd_sc_hd__dfrtp_1 _1904_ (.CLK(clknet_4_15_0_clk),
    .D(_0267_),
    .RESET_B(_0068_),
    .Q(net124));
 sky130_fd_sc_hd__dfrtp_1 _1905_ (.CLK(clknet_4_13_0_clk),
    .D(_0268_),
    .RESET_B(_0069_),
    .Q(net125));
 sky130_fd_sc_hd__dfrtp_1 _1906_ (.CLK(clknet_4_13_0_clk),
    .D(_0269_),
    .RESET_B(_0070_),
    .Q(net126));
 sky130_fd_sc_hd__dfrtp_1 _1907_ (.CLK(clknet_4_12_0_clk),
    .D(_0270_),
    .RESET_B(_0071_),
    .Q(net127));
 sky130_fd_sc_hd__dfrtp_2 _1908_ (.CLK(clknet_4_6_0_clk),
    .D(_0271_),
    .RESET_B(_0072_),
    .Q(\temp_product[32] ));
 sky130_fd_sc_hd__dfrtp_4 _1909_ (.CLK(clknet_4_12_0_clk),
    .D(_0272_),
    .RESET_B(_0073_),
    .Q(\temp_product[33] ));
 sky130_fd_sc_hd__dfrtp_2 _1910_ (.CLK(clknet_4_12_0_clk),
    .D(_0273_),
    .RESET_B(_0074_),
    .Q(\temp_product[34] ));
 sky130_fd_sc_hd__dfrtp_2 _1911_ (.CLK(clknet_4_12_0_clk),
    .D(_0274_),
    .RESET_B(_0075_),
    .Q(\temp_product[35] ));
 sky130_fd_sc_hd__dfrtp_2 _1912_ (.CLK(clknet_4_5_0_clk),
    .D(_0275_),
    .RESET_B(_0076_),
    .Q(\temp_product[36] ));
 sky130_fd_sc_hd__dfrtp_2 _1913_ (.CLK(clknet_4_6_0_clk),
    .D(_0276_),
    .RESET_B(_0077_),
    .Q(\temp_product[37] ));
 sky130_fd_sc_hd__dfrtp_2 _1914_ (.CLK(clknet_4_5_0_clk),
    .D(_0277_),
    .RESET_B(_0078_),
    .Q(\temp_product[38] ));
 sky130_fd_sc_hd__dfrtp_2 _1915_ (.CLK(clknet_4_7_0_clk),
    .D(_0278_),
    .RESET_B(_0079_),
    .Q(\temp_product[39] ));
 sky130_fd_sc_hd__dfrtp_2 _1916_ (.CLK(clknet_4_7_0_clk),
    .D(_0279_),
    .RESET_B(_0080_),
    .Q(\temp_product[40] ));
 sky130_fd_sc_hd__dfrtp_2 _1917_ (.CLK(clknet_4_5_0_clk),
    .D(_0280_),
    .RESET_B(_0081_),
    .Q(\temp_product[41] ));
 sky130_fd_sc_hd__dfrtp_1 _1918_ (.CLK(clknet_4_7_0_clk),
    .D(_0281_),
    .RESET_B(_0082_),
    .Q(\temp_product[42] ));
 sky130_fd_sc_hd__dfrtp_1 _1919_ (.CLK(clknet_4_5_0_clk),
    .D(_0282_),
    .RESET_B(_0083_),
    .Q(\temp_product[43] ));
 sky130_fd_sc_hd__dfrtp_2 _1920_ (.CLK(clknet_4_7_0_clk),
    .D(_0283_),
    .RESET_B(_0084_),
    .Q(\temp_product[44] ));
 sky130_fd_sc_hd__dfrtp_2 _1921_ (.CLK(clknet_4_7_0_clk),
    .D(_0284_),
    .RESET_B(_0085_),
    .Q(\temp_product[45] ));
 sky130_fd_sc_hd__dfrtp_1 _1922_ (.CLK(clknet_4_7_0_clk),
    .D(_0285_),
    .RESET_B(_0086_),
    .Q(\temp_product[46] ));
 sky130_fd_sc_hd__dfrtp_2 _1923_ (.CLK(clknet_4_13_0_clk),
    .D(_0286_),
    .RESET_B(_0087_),
    .Q(\temp_product[47] ));
 sky130_fd_sc_hd__dfrtp_2 _1924_ (.CLK(clknet_4_12_0_clk),
    .D(_0287_),
    .RESET_B(_0088_),
    .Q(\temp_product[48] ));
 sky130_fd_sc_hd__dfrtp_4 _1925_ (.CLK(clknet_4_14_0_clk),
    .D(_0288_),
    .RESET_B(_0089_),
    .Q(\temp_product[49] ));
 sky130_fd_sc_hd__dfrtp_1 _1926_ (.CLK(clknet_4_14_0_clk),
    .D(_0289_),
    .RESET_B(_0090_),
    .Q(\temp_product[50] ));
 sky130_fd_sc_hd__dfrtp_1 _1927_ (.CLK(clknet_4_14_0_clk),
    .D(_0290_),
    .RESET_B(_0091_),
    .Q(\temp_product[51] ));
 sky130_fd_sc_hd__dfrtp_2 _1928_ (.CLK(clknet_4_13_0_clk),
    .D(_0291_),
    .RESET_B(_0092_),
    .Q(\temp_product[52] ));
 sky130_fd_sc_hd__dfrtp_2 _1929_ (.CLK(clknet_4_13_0_clk),
    .D(_0292_),
    .RESET_B(_0093_),
    .Q(\temp_product[53] ));
 sky130_fd_sc_hd__dfrtp_1 _1930_ (.CLK(clknet_4_14_0_clk),
    .D(_0293_),
    .RESET_B(_0094_),
    .Q(\temp_product[54] ));
 sky130_fd_sc_hd__dfrtp_1 _1931_ (.CLK(clknet_4_15_0_clk),
    .D(_0294_),
    .RESET_B(_0095_),
    .Q(\temp_product[55] ));
 sky130_fd_sc_hd__dfrtp_4 _1932_ (.CLK(clknet_4_15_0_clk),
    .D(_0295_),
    .RESET_B(_0096_),
    .Q(\temp_product[56] ));
 sky130_fd_sc_hd__dfrtp_2 _1933_ (.CLK(clknet_4_15_0_clk),
    .D(_0296_),
    .RESET_B(_0097_),
    .Q(\temp_product[57] ));
 sky130_fd_sc_hd__dfrtp_1 _1934_ (.CLK(clknet_4_15_0_clk),
    .D(_0297_),
    .RESET_B(_0098_),
    .Q(\temp_product[58] ));
 sky130_fd_sc_hd__dfrtp_1 _1935_ (.CLK(clknet_4_15_0_clk),
    .D(_0298_),
    .RESET_B(_0099_),
    .Q(\temp_product[59] ));
 sky130_fd_sc_hd__dfrtp_1 _1936_ (.CLK(clknet_4_15_0_clk),
    .D(_0299_),
    .RESET_B(_0100_),
    .Q(\temp_product[60] ));
 sky130_fd_sc_hd__dfrtp_1 _1937_ (.CLK(clknet_4_13_0_clk),
    .D(_0300_),
    .RESET_B(_0101_),
    .Q(\temp_product[61] ));
 sky130_fd_sc_hd__dfrtp_1 _1938_ (.CLK(clknet_4_13_0_clk),
    .D(_0301_),
    .RESET_B(_0102_),
    .Q(\temp_product[62] ));
 sky130_fd_sc_hd__dfrtp_1 _1939_ (.CLK(clknet_4_13_0_clk),
    .D(_0302_),
    .RESET_B(_0103_),
    .Q(\temp_product[63] ));
 sky130_fd_sc_hd__dfrtp_2 _1940_ (.CLK(clknet_4_4_0_clk),
    .D(_0303_),
    .RESET_B(_0104_),
    .Q(\a[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1941_ (.CLK(clknet_4_1_0_clk),
    .D(_0304_),
    .RESET_B(_0105_),
    .Q(\a[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1942_ (.CLK(clknet_4_1_0_clk),
    .D(_0305_),
    .RESET_B(_0106_),
    .Q(\a[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1943_ (.CLK(clknet_4_0_0_clk),
    .D(_0306_),
    .RESET_B(_0107_),
    .Q(\a[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1944_ (.CLK(clknet_4_0_0_clk),
    .D(_0307_),
    .RESET_B(_0108_),
    .Q(\a[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1945_ (.CLK(clknet_4_0_0_clk),
    .D(_0308_),
    .RESET_B(_0109_),
    .Q(\a[5] ));
 sky130_fd_sc_hd__dfrtp_2 _1946_ (.CLK(clknet_4_0_0_clk),
    .D(_0309_),
    .RESET_B(_0110_),
    .Q(\a[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1947_ (.CLK(clknet_4_2_0_clk),
    .D(_0310_),
    .RESET_B(_0111_),
    .Q(\a[7] ));
 sky130_fd_sc_hd__dfrtp_1 _1948_ (.CLK(clknet_4_2_0_clk),
    .D(_0311_),
    .RESET_B(_0112_),
    .Q(\a[8] ));
 sky130_fd_sc_hd__dfrtp_1 _1949_ (.CLK(clknet_4_2_0_clk),
    .D(_0312_),
    .RESET_B(_0113_),
    .Q(\a[9] ));
 sky130_fd_sc_hd__dfrtp_1 _1950_ (.CLK(clknet_4_8_0_clk),
    .D(_0313_),
    .RESET_B(_0114_),
    .Q(\a[10] ));
 sky130_fd_sc_hd__dfrtp_1 _1951_ (.CLK(clknet_4_8_0_clk),
    .D(_0314_),
    .RESET_B(_0115_),
    .Q(\a[11] ));
 sky130_fd_sc_hd__dfrtp_1 _1952_ (.CLK(clknet_4_8_0_clk),
    .D(_0315_),
    .RESET_B(_0116_),
    .Q(\a[12] ));
 sky130_fd_sc_hd__dfrtp_2 _1953_ (.CLK(clknet_4_8_0_clk),
    .D(_0316_),
    .RESET_B(_0117_),
    .Q(\a[13] ));
 sky130_fd_sc_hd__dfrtp_2 _1954_ (.CLK(clknet_4_10_0_clk),
    .D(_0317_),
    .RESET_B(_0118_),
    .Q(\a[14] ));
 sky130_fd_sc_hd__dfrtp_1 _1955_ (.CLK(clknet_4_8_0_clk),
    .D(_0318_),
    .RESET_B(_0119_),
    .Q(\a[15] ));
 sky130_fd_sc_hd__dfrtp_2 _1956_ (.CLK(clknet_4_8_0_clk),
    .D(_0319_),
    .RESET_B(_0120_),
    .Q(\a[16] ));
 sky130_fd_sc_hd__dfrtp_1 _1957_ (.CLK(clknet_4_9_0_clk),
    .D(_0320_),
    .RESET_B(_0121_),
    .Q(\a[17] ));
 sky130_fd_sc_hd__dfrtp_1 _1958_ (.CLK(clknet_4_8_0_clk),
    .D(_0321_),
    .RESET_B(_0122_),
    .Q(\a[18] ));
 sky130_fd_sc_hd__dfrtp_1 _1959_ (.CLK(clknet_4_10_0_clk),
    .D(_0322_),
    .RESET_B(_0123_),
    .Q(\a[19] ));
 sky130_fd_sc_hd__dfrtp_1 _1960_ (.CLK(clknet_4_11_0_clk),
    .D(_0323_),
    .RESET_B(_0124_),
    .Q(\a[20] ));
 sky130_fd_sc_hd__dfrtp_2 _1961_ (.CLK(clknet_4_11_0_clk),
    .D(_0324_),
    .RESET_B(_0125_),
    .Q(\a[21] ));
 sky130_fd_sc_hd__dfrtp_1 _1962_ (.CLK(clknet_4_11_0_clk),
    .D(_0325_),
    .RESET_B(_0126_),
    .Q(\a[22] ));
 sky130_fd_sc_hd__dfrtp_1 _1963_ (.CLK(clknet_4_11_0_clk),
    .D(_0326_),
    .RESET_B(_0127_),
    .Q(\a[23] ));
 sky130_fd_sc_hd__dfrtp_1 _1964_ (.CLK(clknet_4_11_0_clk),
    .D(_0327_),
    .RESET_B(_0128_),
    .Q(\a[24] ));
 sky130_fd_sc_hd__dfrtp_2 _1965_ (.CLK(clknet_4_9_0_clk),
    .D(_0328_),
    .RESET_B(_0129_),
    .Q(\a[25] ));
 sky130_fd_sc_hd__dfrtp_1 _1966_ (.CLK(clknet_4_9_0_clk),
    .D(_0329_),
    .RESET_B(_0130_),
    .Q(\a[26] ));
 sky130_fd_sc_hd__dfrtp_1 _1967_ (.CLK(clknet_4_3_0_clk),
    .D(_0330_),
    .RESET_B(_0131_),
    .Q(\a[27] ));
 sky130_fd_sc_hd__dfrtp_1 _1968_ (.CLK(clknet_4_3_0_clk),
    .D(_0331_),
    .RESET_B(_0132_),
    .Q(\a[28] ));
 sky130_fd_sc_hd__dfrtp_1 _1969_ (.CLK(clknet_4_3_0_clk),
    .D(_0332_),
    .RESET_B(_0133_),
    .Q(\a[29] ));
 sky130_fd_sc_hd__dfrtp_1 _1970_ (.CLK(clknet_4_3_0_clk),
    .D(_0333_),
    .RESET_B(_0134_),
    .Q(\a[30] ));
 sky130_fd_sc_hd__dfrtp_1 _1971_ (.CLK(clknet_4_6_0_clk),
    .D(_0334_),
    .RESET_B(_0135_),
    .Q(\a[31] ));
 sky130_fd_sc_hd__dfrtp_1 _1972_ (.CLK(clknet_4_4_0_clk),
    .D(_0335_),
    .RESET_B(_0136_),
    .Q(\b[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1973_ (.CLK(clknet_4_5_0_clk),
    .D(_0336_),
    .RESET_B(_0137_),
    .Q(\b[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1974_ (.CLK(clknet_4_5_0_clk),
    .D(_0337_),
    .RESET_B(_0138_),
    .Q(\b[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1975_ (.CLK(clknet_4_5_0_clk),
    .D(_0338_),
    .RESET_B(_0139_),
    .Q(\b[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1976_ (.CLK(clknet_4_1_0_clk),
    .D(_0339_),
    .RESET_B(_0140_),
    .Q(\b[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1977_ (.CLK(clknet_4_1_0_clk),
    .D(_0340_),
    .RESET_B(_0141_),
    .Q(\b[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1978_ (.CLK(clknet_4_1_0_clk),
    .D(_0341_),
    .RESET_B(_0142_),
    .Q(\b[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1979_ (.CLK(clknet_4_1_0_clk),
    .D(_0342_),
    .RESET_B(_0143_),
    .Q(\b[7] ));
 sky130_fd_sc_hd__dfrtp_1 _1980_ (.CLK(clknet_4_0_0_clk),
    .D(_0343_),
    .RESET_B(_0144_),
    .Q(\b[8] ));
 sky130_fd_sc_hd__dfrtp_1 _1981_ (.CLK(clknet_4_0_0_clk),
    .D(_0344_),
    .RESET_B(_0145_),
    .Q(\b[9] ));
 sky130_fd_sc_hd__dfrtp_1 _1982_ (.CLK(clknet_4_0_0_clk),
    .D(_0345_),
    .RESET_B(_0146_),
    .Q(\b[10] ));
 sky130_fd_sc_hd__dfrtp_1 _1983_ (.CLK(clknet_4_0_0_clk),
    .D(_0346_),
    .RESET_B(_0147_),
    .Q(\b[11] ));
 sky130_fd_sc_hd__dfrtp_1 _1984_ (.CLK(clknet_4_0_0_clk),
    .D(_0347_),
    .RESET_B(_0148_),
    .Q(\b[12] ));
 sky130_fd_sc_hd__dfrtp_1 _1985_ (.CLK(clknet_4_0_0_clk),
    .D(_0348_),
    .RESET_B(_0149_),
    .Q(\b[13] ));
 sky130_fd_sc_hd__dfrtp_1 _1986_ (.CLK(clknet_4_0_0_clk),
    .D(_0349_),
    .RESET_B(_0150_),
    .Q(\b[14] ));
 sky130_fd_sc_hd__dfrtp_1 _1987_ (.CLK(clknet_4_0_0_clk),
    .D(_0350_),
    .RESET_B(_0151_),
    .Q(\b[15] ));
 sky130_fd_sc_hd__dfrtp_1 _1988_ (.CLK(clknet_4_1_0_clk),
    .D(_0351_),
    .RESET_B(_0152_),
    .Q(\b[16] ));
 sky130_fd_sc_hd__dfrtp_1 _1989_ (.CLK(clknet_4_1_0_clk),
    .D(_0352_),
    .RESET_B(_0153_),
    .Q(\b[17] ));
 sky130_fd_sc_hd__dfrtp_1 _1990_ (.CLK(clknet_4_1_0_clk),
    .D(_0353_),
    .RESET_B(_0154_),
    .Q(\b[18] ));
 sky130_fd_sc_hd__dfrtp_1 _1991_ (.CLK(clknet_4_1_0_clk),
    .D(_0354_),
    .RESET_B(_0155_),
    .Q(\b[19] ));
 sky130_fd_sc_hd__dfrtp_1 _1992_ (.CLK(clknet_4_4_0_clk),
    .D(_0355_),
    .RESET_B(_0156_),
    .Q(\b[20] ));
 sky130_fd_sc_hd__dfrtp_1 _1993_ (.CLK(clknet_4_4_0_clk),
    .D(_0356_),
    .RESET_B(_0157_),
    .Q(\b[21] ));
 sky130_fd_sc_hd__dfrtp_1 _1994_ (.CLK(clknet_4_4_0_clk),
    .D(_0357_),
    .RESET_B(_0158_),
    .Q(\b[22] ));
 sky130_fd_sc_hd__dfrtp_1 _1995_ (.CLK(clknet_4_5_0_clk),
    .D(_0358_),
    .RESET_B(_0159_),
    .Q(\b[23] ));
 sky130_fd_sc_hd__dfrtp_1 _1996_ (.CLK(clknet_4_5_0_clk),
    .D(_0359_),
    .RESET_B(_0160_),
    .Q(\b[24] ));
 sky130_fd_sc_hd__dfrtp_1 _1997_ (.CLK(clknet_4_5_0_clk),
    .D(_0360_),
    .RESET_B(_0161_),
    .Q(\b[25] ));
 sky130_fd_sc_hd__dfrtp_1 _1998_ (.CLK(clknet_4_5_0_clk),
    .D(_0361_),
    .RESET_B(_0162_),
    .Q(\b[26] ));
 sky130_fd_sc_hd__dfrtp_1 _1999_ (.CLK(clknet_4_6_0_clk),
    .D(_0362_),
    .RESET_B(_0163_),
    .Q(\b[27] ));
 sky130_fd_sc_hd__dfrtp_1 _2000_ (.CLK(clknet_4_5_0_clk),
    .D(_0363_),
    .RESET_B(_0164_),
    .Q(\b[28] ));
 sky130_fd_sc_hd__dfrtp_1 _2001_ (.CLK(clknet_4_4_0_clk),
    .D(_0364_),
    .RESET_B(_0165_),
    .Q(\b[29] ));
 sky130_fd_sc_hd__dfrtp_1 _2002_ (.CLK(clknet_4_4_0_clk),
    .D(_0365_),
    .RESET_B(_0166_),
    .Q(\b[30] ));
 sky130_fd_sc_hd__dfrtp_2 _2003_ (.CLK(clknet_4_4_0_clk),
    .D(_0366_),
    .RESET_B(_0167_),
    .Q(\temp_product[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2004_ (.CLK(clknet_4_3_0_clk),
    .D(_0367_),
    .RESET_B(_0168_),
    .Q(\temp_product[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2005_ (.CLK(clknet_4_1_0_clk),
    .D(_0368_),
    .RESET_B(_0169_),
    .Q(\temp_product[2] ));
 sky130_fd_sc_hd__dfrtp_1 _2006_ (.CLK(clknet_4_0_0_clk),
    .D(_0369_),
    .RESET_B(_0170_),
    .Q(\temp_product[3] ));
 sky130_fd_sc_hd__dfrtp_2 _2007_ (.CLK(clknet_4_2_0_clk),
    .D(_0370_),
    .RESET_B(_0171_),
    .Q(\temp_product[4] ));
 sky130_fd_sc_hd__dfrtp_1 _2008_ (.CLK(clknet_4_0_0_clk),
    .D(_0371_),
    .RESET_B(_0172_),
    .Q(\temp_product[5] ));
 sky130_fd_sc_hd__dfrtp_2 _2009_ (.CLK(clknet_4_2_0_clk),
    .D(_0372_),
    .RESET_B(_0173_),
    .Q(\temp_product[6] ));
 sky130_fd_sc_hd__dfrtp_1 _2010_ (.CLK(clknet_4_0_0_clk),
    .D(_0373_),
    .RESET_B(_0174_),
    .Q(\temp_product[7] ));
 sky130_fd_sc_hd__dfrtp_1 _2011_ (.CLK(clknet_4_3_0_clk),
    .D(_0374_),
    .RESET_B(_0175_),
    .Q(\temp_product[8] ));
 sky130_fd_sc_hd__dfrtp_1 _2012_ (.CLK(clknet_4_2_0_clk),
    .D(_0375_),
    .RESET_B(_0176_),
    .Q(\temp_product[9] ));
 sky130_fd_sc_hd__dfrtp_1 _2013_ (.CLK(clknet_4_8_0_clk),
    .D(_0376_),
    .RESET_B(_0177_),
    .Q(\temp_product[10] ));
 sky130_fd_sc_hd__dfrtp_2 _2014_ (.CLK(clknet_4_9_0_clk),
    .D(_0377_),
    .RESET_B(_0178_),
    .Q(\temp_product[11] ));
 sky130_fd_sc_hd__dfrtp_1 _2015_ (.CLK(clknet_4_8_0_clk),
    .D(_0378_),
    .RESET_B(_0179_),
    .Q(\temp_product[12] ));
 sky130_fd_sc_hd__dfrtp_2 _2016_ (.CLK(clknet_4_10_0_clk),
    .D(_0379_),
    .RESET_B(_0180_),
    .Q(\temp_product[13] ));
 sky130_fd_sc_hd__dfrtp_1 _2017_ (.CLK(clknet_4_10_0_clk),
    .D(_0380_),
    .RESET_B(_0181_),
    .Q(\temp_product[14] ));
 sky130_fd_sc_hd__dfrtp_1 _2018_ (.CLK(clknet_4_10_0_clk),
    .D(_0381_),
    .RESET_B(_0182_),
    .Q(\temp_product[15] ));
 sky130_fd_sc_hd__dfrtp_2 _2019_ (.CLK(clknet_4_9_0_clk),
    .D(_0382_),
    .RESET_B(_0183_),
    .Q(\temp_product[16] ));
 sky130_fd_sc_hd__dfrtp_1 _2020_ (.CLK(clknet_4_10_0_clk),
    .D(_0383_),
    .RESET_B(_0184_),
    .Q(\temp_product[17] ));
 sky130_fd_sc_hd__dfrtp_1 _2021_ (.CLK(clknet_4_10_0_clk),
    .D(_0384_),
    .RESET_B(_0185_),
    .Q(\temp_product[18] ));
 sky130_fd_sc_hd__dfrtp_1 _2022_ (.CLK(clknet_4_10_0_clk),
    .D(_0385_),
    .RESET_B(_0186_),
    .Q(\temp_product[19] ));
 sky130_fd_sc_hd__dfrtp_1 _2023_ (.CLK(clknet_4_10_0_clk),
    .D(_0386_),
    .RESET_B(_0187_),
    .Q(\temp_product[20] ));
 sky130_fd_sc_hd__dfrtp_2 _2024_ (.CLK(clknet_4_11_0_clk),
    .D(_0387_),
    .RESET_B(_0188_),
    .Q(\temp_product[21] ));
 sky130_fd_sc_hd__dfrtp_1 _2025_ (.CLK(clknet_4_11_0_clk),
    .D(_0388_),
    .RESET_B(_0189_),
    .Q(\temp_product[22] ));
 sky130_fd_sc_hd__dfrtp_1 _2026_ (.CLK(clknet_4_9_0_clk),
    .D(_0389_),
    .RESET_B(_0190_),
    .Q(\temp_product[23] ));
 sky130_fd_sc_hd__dfrtp_1 _2027_ (.CLK(clknet_4_9_0_clk),
    .D(_0390_),
    .RESET_B(_0191_),
    .Q(\temp_product[24] ));
 sky130_fd_sc_hd__dfrtp_2 _2028_ (.CLK(clknet_4_9_0_clk),
    .D(_0391_),
    .RESET_B(_0192_),
    .Q(\temp_product[25] ));
 sky130_fd_sc_hd__dfrtp_1 _2029_ (.CLK(clknet_4_9_0_clk),
    .D(_0392_),
    .RESET_B(_0193_),
    .Q(\temp_product[26] ));
 sky130_fd_sc_hd__dfrtp_1 _2030_ (.CLK(clknet_4_3_0_clk),
    .D(_0393_),
    .RESET_B(_0194_),
    .Q(\temp_product[27] ));
 sky130_fd_sc_hd__dfrtp_1 _2031_ (.CLK(clknet_4_3_0_clk),
    .D(_0394_),
    .RESET_B(_0195_),
    .Q(\temp_product[28] ));
 sky130_fd_sc_hd__dfrtp_1 _2032_ (.CLK(clknet_4_3_0_clk),
    .D(_0395_),
    .RESET_B(_0196_),
    .Q(\temp_product[29] ));
 sky130_fd_sc_hd__dfrtp_2 _2033_ (.CLK(clknet_4_6_0_clk),
    .D(_0396_),
    .RESET_B(_0197_),
    .Q(\temp_product[30] ));
 sky130_fd_sc_hd__dfrtp_1 _2034_ (.CLK(clknet_4_3_0_clk),
    .D(_0397_),
    .RESET_B(_0198_),
    .Q(\temp_product[31] ));
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(multiplicand[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(multiplicand[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(multiplicand[11]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(multiplicand[12]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(multiplicand[13]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(multiplicand[14]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(multiplicand[15]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(multiplicand[16]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(multiplicand[17]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(multiplicand[18]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(multiplicand[19]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(multiplicand[1]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(multiplicand[20]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(multiplicand[21]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(multiplicand[22]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(multiplicand[23]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(multiplicand[24]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(multiplicand[25]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(multiplicand[26]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(multiplicand[27]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(multiplicand[28]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(multiplicand[29]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(multiplicand[2]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(multiplicand[30]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_2 input25 (.A(multiplicand[31]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(multiplicand[3]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(multiplicand[4]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(multiplicand[5]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(multiplicand[6]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(multiplicand[7]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(multiplicand[8]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(multiplicand[9]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(multiplier[0]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(multiplier[10]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(multiplier[11]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(multiplier[12]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(multiplier[13]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 input38 (.A(multiplier[14]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 input39 (.A(multiplier[15]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(multiplier[16]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 input41 (.A(multiplier[17]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 input42 (.A(multiplier[18]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 input43 (.A(multiplier[19]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(multiplier[1]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(multiplier[20]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_1 input46 (.A(multiplier[21]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_1 input47 (.A(multiplier[22]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_1 input48 (.A(multiplier[23]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_1 input49 (.A(multiplier[24]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_1 input50 (.A(multiplier[25]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 input51 (.A(multiplier[26]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_1 input52 (.A(multiplier[27]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 input53 (.A(multiplier[28]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 input54 (.A(multiplier[29]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_1 input55 (.A(multiplier[2]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_1 input56 (.A(multiplier[30]),
    .X(net56));
 sky130_fd_sc_hd__buf_1 input57 (.A(multiplier[31]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_1 input58 (.A(multiplier[3]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 input59 (.A(multiplier[4]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_1 input60 (.A(multiplier[5]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_1 input61 (.A(multiplier[6]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 input62 (.A(multiplier[7]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_1 input63 (.A(multiplier[8]),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_1 input64 (.A(multiplier[9]),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_1 input65 (.A(rst),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_1 input66 (.A(start),
    .X(net66));
 sky130_fd_sc_hd__buf_2 output67 (.A(net67),
    .X(done));
 sky130_fd_sc_hd__buf_2 output68 (.A(net68),
    .X(product[0]));
 sky130_fd_sc_hd__buf_2 output69 (.A(net69),
    .X(product[10]));
 sky130_fd_sc_hd__buf_2 output70 (.A(net70),
    .X(product[11]));
 sky130_fd_sc_hd__buf_2 output71 (.A(net71),
    .X(product[12]));
 sky130_fd_sc_hd__buf_2 output72 (.A(net72),
    .X(product[13]));
 sky130_fd_sc_hd__buf_2 output73 (.A(net73),
    .X(product[14]));
 sky130_fd_sc_hd__buf_2 output74 (.A(net74),
    .X(product[15]));
 sky130_fd_sc_hd__buf_2 output75 (.A(net75),
    .X(product[16]));
 sky130_fd_sc_hd__buf_2 output76 (.A(net76),
    .X(product[17]));
 sky130_fd_sc_hd__buf_2 output77 (.A(net77),
    .X(product[18]));
 sky130_fd_sc_hd__buf_2 output78 (.A(net78),
    .X(product[19]));
 sky130_fd_sc_hd__buf_2 output79 (.A(net79),
    .X(product[1]));
 sky130_fd_sc_hd__buf_2 output80 (.A(net80),
    .X(product[20]));
 sky130_fd_sc_hd__buf_2 output81 (.A(net81),
    .X(product[21]));
 sky130_fd_sc_hd__buf_2 output82 (.A(net82),
    .X(product[22]));
 sky130_fd_sc_hd__buf_2 output83 (.A(net83),
    .X(product[23]));
 sky130_fd_sc_hd__buf_2 output84 (.A(net84),
    .X(product[24]));
 sky130_fd_sc_hd__buf_2 output85 (.A(net85),
    .X(product[25]));
 sky130_fd_sc_hd__buf_2 output86 (.A(net86),
    .X(product[26]));
 sky130_fd_sc_hd__buf_2 output87 (.A(net87),
    .X(product[27]));
 sky130_fd_sc_hd__buf_2 output88 (.A(net88),
    .X(product[28]));
 sky130_fd_sc_hd__buf_2 output89 (.A(net89),
    .X(product[29]));
 sky130_fd_sc_hd__buf_2 output90 (.A(net90),
    .X(product[2]));
 sky130_fd_sc_hd__buf_2 output91 (.A(net91),
    .X(product[30]));
 sky130_fd_sc_hd__buf_2 output92 (.A(net92),
    .X(product[31]));
 sky130_fd_sc_hd__buf_2 output93 (.A(net93),
    .X(product[32]));
 sky130_fd_sc_hd__buf_2 output94 (.A(net94),
    .X(product[33]));
 sky130_fd_sc_hd__buf_2 output95 (.A(net95),
    .X(product[34]));
 sky130_fd_sc_hd__buf_2 output96 (.A(net96),
    .X(product[35]));
 sky130_fd_sc_hd__buf_2 output97 (.A(net97),
    .X(product[36]));
 sky130_fd_sc_hd__buf_2 output98 (.A(net98),
    .X(product[37]));
 sky130_fd_sc_hd__buf_2 output99 (.A(net99),
    .X(product[38]));
 sky130_fd_sc_hd__buf_2 output100 (.A(net100),
    .X(product[39]));
 sky130_fd_sc_hd__buf_2 output101 (.A(net101),
    .X(product[3]));
 sky130_fd_sc_hd__buf_2 output102 (.A(net102),
    .X(product[40]));
 sky130_fd_sc_hd__buf_2 output103 (.A(net103),
    .X(product[41]));
 sky130_fd_sc_hd__buf_2 output104 (.A(net104),
    .X(product[42]));
 sky130_fd_sc_hd__buf_2 output105 (.A(net105),
    .X(product[43]));
 sky130_fd_sc_hd__buf_2 output106 (.A(net106),
    .X(product[44]));
 sky130_fd_sc_hd__buf_2 output107 (.A(net107),
    .X(product[45]));
 sky130_fd_sc_hd__buf_2 output108 (.A(net108),
    .X(product[46]));
 sky130_fd_sc_hd__buf_2 output109 (.A(net109),
    .X(product[47]));
 sky130_fd_sc_hd__buf_2 output110 (.A(net110),
    .X(product[48]));
 sky130_fd_sc_hd__buf_2 output111 (.A(net111),
    .X(product[49]));
 sky130_fd_sc_hd__buf_2 output112 (.A(net112),
    .X(product[4]));
 sky130_fd_sc_hd__buf_2 output113 (.A(net113),
    .X(product[50]));
 sky130_fd_sc_hd__buf_2 output114 (.A(net114),
    .X(product[51]));
 sky130_fd_sc_hd__buf_2 output115 (.A(net115),
    .X(product[52]));
 sky130_fd_sc_hd__buf_2 output116 (.A(net116),
    .X(product[53]));
 sky130_fd_sc_hd__buf_2 output117 (.A(net117),
    .X(product[54]));
 sky130_fd_sc_hd__buf_2 output118 (.A(net118),
    .X(product[55]));
 sky130_fd_sc_hd__buf_2 output119 (.A(net119),
    .X(product[56]));
 sky130_fd_sc_hd__buf_2 output120 (.A(net120),
    .X(product[57]));
 sky130_fd_sc_hd__buf_2 output121 (.A(net121),
    .X(product[58]));
 sky130_fd_sc_hd__buf_2 output122 (.A(net122),
    .X(product[59]));
 sky130_fd_sc_hd__buf_2 output123 (.A(net123),
    .X(product[5]));
 sky130_fd_sc_hd__buf_2 output124 (.A(net124),
    .X(product[60]));
 sky130_fd_sc_hd__buf_2 output125 (.A(net125),
    .X(product[61]));
 sky130_fd_sc_hd__buf_2 output126 (.A(net126),
    .X(product[62]));
 sky130_fd_sc_hd__buf_2 output127 (.A(net127),
    .X(product[63]));
 sky130_fd_sc_hd__buf_2 output128 (.A(net128),
    .X(product[6]));
 sky130_fd_sc_hd__buf_2 output129 (.A(net129),
    .X(product[7]));
 sky130_fd_sc_hd__buf_2 output130 (.A(net130),
    .X(product[8]));
 sky130_fd_sc_hd__buf_2 output131 (.A(net131),
    .X(product[9]));
 sky130_fd_sc_hd__buf_2 fanout132 (.A(_0676_),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_2 fanout133 (.A(_0676_),
    .X(net133));
 sky130_fd_sc_hd__buf_2 fanout134 (.A(_0676_),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_2 fanout135 (.A(_0676_),
    .X(net135));
 sky130_fd_sc_hd__buf_2 fanout136 (.A(net137),
    .X(net136));
 sky130_fd_sc_hd__clkbuf_4 fanout137 (.A(_0409_),
    .X(net137));
 sky130_fd_sc_hd__buf_2 fanout138 (.A(net140),
    .X(net138));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout139 (.A(net140),
    .X(net139));
 sky130_fd_sc_hd__clkbuf_2 fanout140 (.A(_0409_),
    .X(net140));
 sky130_fd_sc_hd__buf_2 fanout141 (.A(net143),
    .X(net141));
 sky130_fd_sc_hd__buf_2 fanout142 (.A(net143),
    .X(net142));
 sky130_fd_sc_hd__clkbuf_2 fanout143 (.A(_0409_),
    .X(net143));
 sky130_fd_sc_hd__buf_2 fanout144 (.A(net147),
    .X(net144));
 sky130_fd_sc_hd__buf_2 fanout145 (.A(net147),
    .X(net145));
 sky130_fd_sc_hd__clkbuf_2 fanout146 (.A(net147),
    .X(net146));
 sky130_fd_sc_hd__clkbuf_2 fanout147 (.A(_0798_),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_4 fanout148 (.A(net151),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_4 fanout149 (.A(net150),
    .X(net149));
 sky130_fd_sc_hd__clkbuf_4 fanout150 (.A(net151),
    .X(net150));
 sky130_fd_sc_hd__clkbuf_2 fanout151 (.A(_0798_),
    .X(net151));
 sky130_fd_sc_hd__clkbuf_4 fanout152 (.A(_0675_),
    .X(net152));
 sky130_fd_sc_hd__clkbuf_2 fanout153 (.A(_0675_),
    .X(net153));
 sky130_fd_sc_hd__buf_2 fanout154 (.A(net155),
    .X(net154));
 sky130_fd_sc_hd__buf_2 fanout155 (.A(_0675_),
    .X(net155));
 sky130_fd_sc_hd__buf_2 fanout156 (.A(net157),
    .X(net156));
 sky130_fd_sc_hd__buf_2 fanout157 (.A(net158),
    .X(net157));
 sky130_fd_sc_hd__clkbuf_2 fanout158 (.A(net161),
    .X(net158));
 sky130_fd_sc_hd__buf_2 fanout159 (.A(net161),
    .X(net159));
 sky130_fd_sc_hd__clkbuf_2 fanout160 (.A(net161),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_2 fanout161 (.A(_0673_),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_4 fanout162 (.A(net164),
    .X(net162));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout163 (.A(net164),
    .X(net163));
 sky130_fd_sc_hd__clkbuf_2 fanout164 (.A(_0673_),
    .X(net164));
 sky130_fd_sc_hd__clkbuf_4 fanout165 (.A(net167),
    .X(net165));
 sky130_fd_sc_hd__clkbuf_4 fanout166 (.A(net167),
    .X(net166));
 sky130_fd_sc_hd__buf_4 fanout167 (.A(_0672_),
    .X(net167));
 sky130_fd_sc_hd__clkbuf_4 fanout168 (.A(net172),
    .X(net168));
 sky130_fd_sc_hd__buf_2 fanout169 (.A(net172),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_2 fanout170 (.A(net172),
    .X(net170));
 sky130_fd_sc_hd__buf_2 fanout171 (.A(net172),
    .X(net171));
 sky130_fd_sc_hd__clkbuf_4 fanout172 (.A(_0672_),
    .X(net172));
 sky130_fd_sc_hd__buf_2 fanout173 (.A(net174),
    .X(net173));
 sky130_fd_sc_hd__buf_2 fanout174 (.A(net175),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_2 fanout175 (.A(net178),
    .X(net175));
 sky130_fd_sc_hd__buf_2 fanout176 (.A(net178),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_2 fanout177 (.A(net178),
    .X(net177));
 sky130_fd_sc_hd__clkbuf_2 fanout178 (.A(_0671_),
    .X(net178));
 sky130_fd_sc_hd__clkbuf_4 fanout179 (.A(net181),
    .X(net179));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout180 (.A(net181),
    .X(net180));
 sky130_fd_sc_hd__clkbuf_2 fanout181 (.A(_0671_),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_4 fanout182 (.A(_0670_),
    .X(net182));
 sky130_fd_sc_hd__buf_2 fanout183 (.A(net185),
    .X(net183));
 sky130_fd_sc_hd__clkbuf_2 fanout184 (.A(net185),
    .X(net184));
 sky130_fd_sc_hd__buf_2 fanout185 (.A(_0669_),
    .X(net185));
 sky130_fd_sc_hd__clkbuf_1 max_cap186 (.A(_0501_),
    .X(net186));
 sky130_fd_sc_hd__buf_2 fanout187 (.A(net191),
    .X(net187));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout188 (.A(net191),
    .X(net188));
 sky130_fd_sc_hd__buf_2 fanout189 (.A(net191),
    .X(net189));
 sky130_fd_sc_hd__clkbuf_2 fanout190 (.A(net191),
    .X(net190));
 sky130_fd_sc_hd__buf_2 fanout191 (.A(\a[31] ),
    .X(net191));
 sky130_fd_sc_hd__buf_2 fanout192 (.A(net193),
    .X(net192));
 sky130_fd_sc_hd__buf_2 fanout193 (.A(net194),
    .X(net193));
 sky130_fd_sc_hd__clkbuf_2 fanout194 (.A(net195),
    .X(net194));
 sky130_fd_sc_hd__buf_2 fanout195 (.A(\a[31] ),
    .X(net195));
 sky130_fd_sc_hd__clkbuf_2 fanout196 (.A(net198),
    .X(net196));
 sky130_fd_sc_hd__buf_1 fanout197 (.A(net198),
    .X(net197));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout198 (.A(net199),
    .X(net198));
 sky130_fd_sc_hd__clkbuf_2 fanout199 (.A(net205),
    .X(net199));
 sky130_fd_sc_hd__clkbuf_2 fanout200 (.A(net201),
    .X(net200));
 sky130_fd_sc_hd__buf_2 fanout201 (.A(net205),
    .X(net201));
 sky130_fd_sc_hd__buf_2 fanout202 (.A(net203),
    .X(net202));
 sky130_fd_sc_hd__clkbuf_2 fanout203 (.A(net204),
    .X(net203));
 sky130_fd_sc_hd__clkbuf_2 fanout204 (.A(net205),
    .X(net204));
 sky130_fd_sc_hd__buf_2 fanout205 (.A(net66),
    .X(net205));
 sky130_fd_sc_hd__buf_4 fanout206 (.A(net213),
    .X(net206));
 sky130_fd_sc_hd__clkbuf_4 fanout207 (.A(net213),
    .X(net207));
 sky130_fd_sc_hd__buf_4 fanout208 (.A(net213),
    .X(net208));
 sky130_fd_sc_hd__buf_2 fanout209 (.A(net213),
    .X(net209));
 sky130_fd_sc_hd__buf_4 fanout210 (.A(net212),
    .X(net210));
 sky130_fd_sc_hd__clkbuf_4 fanout211 (.A(net212),
    .X(net211));
 sky130_fd_sc_hd__clkbuf_4 fanout212 (.A(net213),
    .X(net212));
 sky130_fd_sc_hd__clkbuf_2 fanout213 (.A(net234),
    .X(net213));
 sky130_fd_sc_hd__buf_4 fanout214 (.A(net220),
    .X(net214));
 sky130_fd_sc_hd__buf_2 fanout215 (.A(net220),
    .X(net215));
 sky130_fd_sc_hd__buf_4 fanout216 (.A(net220),
    .X(net216));
 sky130_fd_sc_hd__buf_2 fanout217 (.A(net220),
    .X(net217));
 sky130_fd_sc_hd__buf_4 fanout218 (.A(net219),
    .X(net218));
 sky130_fd_sc_hd__buf_4 fanout219 (.A(net220),
    .X(net219));
 sky130_fd_sc_hd__buf_2 fanout220 (.A(net234),
    .X(net220));
 sky130_fd_sc_hd__buf_4 fanout221 (.A(net223),
    .X(net221));
 sky130_fd_sc_hd__clkbuf_4 fanout222 (.A(net223),
    .X(net222));
 sky130_fd_sc_hd__clkbuf_4 fanout223 (.A(net226),
    .X(net223));
 sky130_fd_sc_hd__buf_4 fanout224 (.A(net225),
    .X(net224));
 sky130_fd_sc_hd__buf_4 fanout225 (.A(net226),
    .X(net225));
 sky130_fd_sc_hd__buf_2 fanout226 (.A(net234),
    .X(net226));
 sky130_fd_sc_hd__buf_4 fanout227 (.A(net229),
    .X(net227));
 sky130_fd_sc_hd__clkbuf_2 fanout228 (.A(net229),
    .X(net228));
 sky130_fd_sc_hd__buf_2 fanout229 (.A(net234),
    .X(net229));
 sky130_fd_sc_hd__buf_4 fanout230 (.A(net231),
    .X(net230));
 sky130_fd_sc_hd__buf_2 fanout231 (.A(net233),
    .X(net231));
 sky130_fd_sc_hd__buf_4 fanout232 (.A(net233),
    .X(net232));
 sky130_fd_sc_hd__buf_2 fanout233 (.A(net234),
    .X(net233));
 sky130_fd_sc_hd__clkbuf_2 fanout234 (.A(net65),
    .X(net234));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload0 (.A(clknet_4_0_0_clk));
 sky130_fd_sc_hd__bufinv_16 clkload1 (.A(clknet_4_1_0_clk));
 sky130_fd_sc_hd__bufinv_16 clkload2 (.A(clknet_4_2_0_clk));
 sky130_fd_sc_hd__inv_6 clkload3 (.A(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload4 (.A(clknet_4_4_0_clk));
 sky130_fd_sc_hd__inv_8 clkload5 (.A(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkinv_4 clkload6 (.A(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload7 (.A(clknet_4_8_0_clk));
 sky130_fd_sc_hd__inv_8 clkload8 (.A(clknet_4_9_0_clk));
 sky130_fd_sc_hd__bufinv_16 clkload9 (.A(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkinv_4 clkload10 (.A(clknet_4_11_0_clk));
 sky130_fd_sc_hd__inv_8 clkload11 (.A(clknet_4_12_0_clk));
 sky130_fd_sc_hd__inv_6 clkload12 (.A(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkinv_4 clkload13 (.A(clknet_4_14_0_clk));
 sky130_fd_sc_hd__bufinv_16 clkload14 (.A(clknet_4_15_0_clk));
endmodule
