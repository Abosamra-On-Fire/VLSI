module multiplier_r (A,
    B,
    P);
 input [31:0] A;
 input [31:0] B;
 output [63:0] P;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;

 sky130_fd_sc_hd__and4_1 _05307_ (.A(net235),
    .B(net227),
    .C(net598),
    .D(net624),
    .X(_00287_));
 sky130_fd_sc_hd__nand4_1 _05308_ (.A(net434),
    .B(net478),
    .C(net341),
    .D(net485),
    .Y(_00298_));
 sky130_fd_sc_hd__a22o_1 _05309_ (.A1(net434),
    .A2(net478),
    .B1(net341),
    .B2(net485),
    .X(_00309_));
 sky130_fd_sc_hd__and2_1 _05310_ (.A(net255),
    .B(net494),
    .X(_00320_));
 sky130_fd_sc_hd__nand3_1 _05311_ (.A(_00298_),
    .B(_00309_),
    .C(_00320_),
    .Y(_00331_));
 sky130_fd_sc_hd__a21o_1 _05312_ (.A1(_00298_),
    .A2(_00309_),
    .B1(_00320_),
    .X(_00342_));
 sky130_fd_sc_hd__and4_1 _05313_ (.A(net434),
    .B(net341),
    .C(net485),
    .D(net494),
    .X(_00353_));
 sky130_fd_sc_hd__nand2_1 _05314_ (.A(net255),
    .B(net514),
    .Y(_00364_));
 sky130_fd_sc_hd__a22oi_2 _05315_ (.A1(net434),
    .A2(net485),
    .B1(net494),
    .B2(net341),
    .Y(_00374_));
 sky130_fd_sc_hd__or3_1 _05316_ (.A(_00353_),
    .B(_00364_),
    .C(_00374_),
    .X(_00385_));
 sky130_fd_sc_hd__o21bai_1 _05317_ (.A1(_00364_),
    .A2(_00374_),
    .B1_N(_00353_),
    .Y(_00396_));
 sky130_fd_sc_hd__nand3_1 _05318_ (.A(_00331_),
    .B(_00342_),
    .C(_00396_),
    .Y(_00407_));
 sky130_fd_sc_hd__a21o_1 _05319_ (.A1(_00331_),
    .A2(_00342_),
    .B1(_00396_),
    .X(_00418_));
 sky130_fd_sc_hd__and4_1 _05320_ (.A(net514),
    .B(net235),
    .C(net227),
    .D(net598),
    .X(_00429_));
 sky130_fd_sc_hd__a22oi_1 _05321_ (.A1(net514),
    .A2(net235),
    .B1(net227),
    .B2(net598),
    .Y(_00440_));
 sky130_fd_sc_hd__or2_1 _05322_ (.A(_00429_),
    .B(_00440_),
    .X(_00451_));
 sky130_fd_sc_hd__nand2_1 _05323_ (.A(net219),
    .B(net624),
    .Y(_00462_));
 sky130_fd_sc_hd__xor2_1 _05324_ (.A(_00451_),
    .B(_00462_),
    .X(_00473_));
 sky130_fd_sc_hd__nand3_1 _05325_ (.A(_00407_),
    .B(_00418_),
    .C(_00473_),
    .Y(_00484_));
 sky130_fd_sc_hd__a21o_1 _05326_ (.A1(_00407_),
    .A2(_00418_),
    .B1(_00473_),
    .X(_00495_));
 sky130_fd_sc_hd__o21ai_1 _05327_ (.A1(_00353_),
    .A2(_00374_),
    .B1(_00364_),
    .Y(_00505_));
 sky130_fd_sc_hd__and4_1 _05328_ (.A(net434),
    .B(net341),
    .C(net494),
    .D(net514),
    .X(_00516_));
 sky130_fd_sc_hd__nand2_1 _05329_ (.A(net255),
    .B(net598),
    .Y(_00527_));
 sky130_fd_sc_hd__a22oi_1 _05330_ (.A1(net434),
    .A2(net494),
    .B1(net514),
    .B2(net341),
    .Y(_00538_));
 sky130_fd_sc_hd__nor2_1 _05331_ (.A(_00516_),
    .B(_00538_),
    .Y(_00549_));
 sky130_fd_sc_hd__o21bai_1 _05332_ (.A1(_00527_),
    .A2(_00538_),
    .B1_N(_00516_),
    .Y(_00560_));
 sky130_fd_sc_hd__and3_1 _05333_ (.A(_00385_),
    .B(_00505_),
    .C(_00560_),
    .X(_00571_));
 sky130_fd_sc_hd__a22oi_1 _05334_ (.A1(net235),
    .A2(net598),
    .B1(net624),
    .B2(net227),
    .Y(_00582_));
 sky130_fd_sc_hd__nor2_1 _05335_ (.A(_00287_),
    .B(_00582_),
    .Y(_00593_));
 sky130_fd_sc_hd__a21o_1 _05336_ (.A1(_00385_),
    .A2(_00505_),
    .B1(_00560_),
    .X(_00604_));
 sky130_fd_sc_hd__nand2b_1 _05337_ (.A_N(_00571_),
    .B(_00604_),
    .Y(_00615_));
 sky130_fd_sc_hd__a21o_1 _05338_ (.A1(_00593_),
    .A2(_00604_),
    .B1(_00571_),
    .X(_00626_));
 sky130_fd_sc_hd__and3_1 _05339_ (.A(_00484_),
    .B(_00495_),
    .C(_00626_),
    .X(_00636_));
 sky130_fd_sc_hd__a21oi_1 _05340_ (.A1(_00484_),
    .A2(_00495_),
    .B1(_00626_),
    .Y(_00647_));
 sky130_fd_sc_hd__nor2_1 _05341_ (.A(_00636_),
    .B(_00647_),
    .Y(_00658_));
 sky130_fd_sc_hd__xnor2_1 _05342_ (.A(_00287_),
    .B(_00658_),
    .Y(_00669_));
 sky130_fd_sc_hd__xnor2_1 _05343_ (.A(_00593_),
    .B(_00615_),
    .Y(_00680_));
 sky130_fd_sc_hd__xnor2_1 _05344_ (.A(_00527_),
    .B(_00549_),
    .Y(_00691_));
 sky130_fd_sc_hd__and4_1 _05345_ (.A(net434),
    .B(net341),
    .C(net514),
    .D(net598),
    .X(_00702_));
 sky130_fd_sc_hd__a22oi_1 _05346_ (.A1(net434),
    .A2(net514),
    .B1(net598),
    .B2(net341),
    .Y(_00713_));
 sky130_fd_sc_hd__and4bb_1 _05347_ (.A_N(_00702_),
    .B_N(_00713_),
    .C(net255),
    .D(net627),
    .X(_00724_));
 sky130_fd_sc_hd__nor2_1 _05348_ (.A(_00702_),
    .B(_00724_),
    .Y(_00735_));
 sky130_fd_sc_hd__and2b_1 _05349_ (.A_N(_00735_),
    .B(_00691_),
    .X(_00746_));
 sky130_fd_sc_hd__xnor2_1 _05350_ (.A(_00691_),
    .B(_00735_),
    .Y(_00757_));
 sky130_fd_sc_hd__and3_1 _05351_ (.A(net235),
    .B(net624),
    .C(_00757_),
    .X(_00768_));
 sky130_fd_sc_hd__o21ai_2 _05352_ (.A1(_00746_),
    .A2(_00768_),
    .B1(_00680_),
    .Y(_00778_));
 sky130_fd_sc_hd__or3_1 _05353_ (.A(_00680_),
    .B(_00746_),
    .C(_00768_),
    .X(_00789_));
 sky130_fd_sc_hd__and2_1 _05354_ (.A(_00778_),
    .B(_00789_),
    .X(_00800_));
 sky130_fd_sc_hd__a21oi_1 _05355_ (.A1(net235),
    .A2(net624),
    .B1(_00757_),
    .Y(_00811_));
 sky130_fd_sc_hd__nor2_1 _05356_ (.A(_00768_),
    .B(_00811_),
    .Y(_00822_));
 sky130_fd_sc_hd__o2bb2a_1 _05357_ (.A1_N(net255),
    .A2_N(net627),
    .B1(_00702_),
    .B2(_00713_),
    .X(_00833_));
 sky130_fd_sc_hd__nor2_1 _05358_ (.A(_00724_),
    .B(_00833_),
    .Y(_00844_));
 sky130_fd_sc_hd__and2_1 _05359_ (.A(net434),
    .B(net627),
    .X(net65));
 sky130_fd_sc_hd__and3_1 _05360_ (.A(net341),
    .B(net598),
    .C(net65),
    .X(_00865_));
 sky130_fd_sc_hd__and2_1 _05361_ (.A(_00844_),
    .B(_00865_),
    .X(_00876_));
 sky130_fd_sc_hd__and2_1 _05362_ (.A(_00822_),
    .B(_00876_),
    .X(_00887_));
 sky130_fd_sc_hd__nand2_1 _05363_ (.A(_00800_),
    .B(_00887_),
    .Y(_00898_));
 sky130_fd_sc_hd__nand2_1 _05364_ (.A(_00778_),
    .B(_00898_),
    .Y(_00909_));
 sky130_fd_sc_hd__and3_1 _05365_ (.A(_00669_),
    .B(_00778_),
    .C(_00898_),
    .X(_00919_));
 sky130_fd_sc_hd__a21oi_1 _05366_ (.A1(_00778_),
    .A2(_00898_),
    .B1(_00669_),
    .Y(_00930_));
 sky130_fd_sc_hd__nor2_1 _05367_ (.A(_00919_),
    .B(_00930_),
    .Y(net120));
 sky130_fd_sc_hd__and4_1 _05368_ (.A(net435),
    .B(net478),
    .C(net342),
    .D(net470),
    .X(_00951_));
 sky130_fd_sc_hd__a22oi_2 _05369_ (.A1(net478),
    .A2(net342),
    .B1(net470),
    .B2(net435),
    .Y(_00962_));
 sky130_fd_sc_hd__nand2_1 _05370_ (.A(net485),
    .B(net255),
    .Y(_00973_));
 sky130_fd_sc_hd__or3_1 _05371_ (.A(_00951_),
    .B(_00962_),
    .C(_00973_),
    .X(_00984_));
 sky130_fd_sc_hd__o21ai_1 _05372_ (.A1(_00951_),
    .A2(_00962_),
    .B1(_00973_),
    .Y(_00995_));
 sky130_fd_sc_hd__a21bo_1 _05373_ (.A1(_00309_),
    .A2(_00320_),
    .B1_N(_00298_),
    .X(_01006_));
 sky130_fd_sc_hd__nand3_1 _05374_ (.A(_00984_),
    .B(_00995_),
    .C(_01006_),
    .Y(_01017_));
 sky130_fd_sc_hd__a21o_1 _05375_ (.A1(_00984_),
    .A2(_00995_),
    .B1(_01006_),
    .X(_01028_));
 sky130_fd_sc_hd__and4_1 _05376_ (.A(net494),
    .B(net514),
    .C(net235),
    .D(net227),
    .X(_01039_));
 sky130_fd_sc_hd__a22oi_1 _05377_ (.A1(net493),
    .A2(net235),
    .B1(net227),
    .B2(net514),
    .Y(_01050_));
 sky130_fd_sc_hd__nor2_1 _05378_ (.A(_01039_),
    .B(_01050_),
    .Y(_01061_));
 sky130_fd_sc_hd__nand2_1 _05379_ (.A(net598),
    .B(net219),
    .Y(_01071_));
 sky130_fd_sc_hd__xnor2_1 _05380_ (.A(_01061_),
    .B(_01071_),
    .Y(_01082_));
 sky130_fd_sc_hd__nand3_1 _05381_ (.A(_01017_),
    .B(_01028_),
    .C(_01082_),
    .Y(_01093_));
 sky130_fd_sc_hd__a21o_1 _05382_ (.A1(_01017_),
    .A2(_01028_),
    .B1(_01082_),
    .X(_01104_));
 sky130_fd_sc_hd__a21bo_1 _05383_ (.A1(_00418_),
    .A2(_00473_),
    .B1_N(_00407_),
    .X(_01115_));
 sky130_fd_sc_hd__and3_1 _05384_ (.A(_01093_),
    .B(_01104_),
    .C(_01115_),
    .X(_01126_));
 sky130_fd_sc_hd__nand3_1 _05385_ (.A(_01093_),
    .B(_01104_),
    .C(_01115_),
    .Y(_01137_));
 sky130_fd_sc_hd__a21o_1 _05386_ (.A1(_01093_),
    .A2(_01104_),
    .B1(_01115_),
    .X(_01148_));
 sky130_fd_sc_hd__o21bai_1 _05387_ (.A1(_00440_),
    .A2(_00462_),
    .B1_N(_00429_),
    .Y(_01159_));
 sky130_fd_sc_hd__nand2_1 _05388_ (.A(net624),
    .B(net207),
    .Y(_01170_));
 sky130_fd_sc_hd__and3_1 _05389_ (.A(net624),
    .B(net207),
    .C(_01159_),
    .X(_01181_));
 sky130_fd_sc_hd__xnor2_1 _05390_ (.A(_01159_),
    .B(_01170_),
    .Y(_01192_));
 sky130_fd_sc_hd__and3_1 _05391_ (.A(_01137_),
    .B(_01148_),
    .C(_01192_),
    .X(_01203_));
 sky130_fd_sc_hd__a21oi_1 _05392_ (.A1(_01137_),
    .A2(_01148_),
    .B1(_01192_),
    .Y(_01214_));
 sky130_fd_sc_hd__nor2_1 _05393_ (.A(_01203_),
    .B(_01214_),
    .Y(_01224_));
 sky130_fd_sc_hd__a21o_1 _05394_ (.A1(_00287_),
    .A2(_00658_),
    .B1(_00636_),
    .X(_01235_));
 sky130_fd_sc_hd__and2_1 _05395_ (.A(_01224_),
    .B(_01235_),
    .X(_01246_));
 sky130_fd_sc_hd__xnor2_1 _05396_ (.A(_01224_),
    .B(_01235_),
    .Y(_01257_));
 sky130_fd_sc_hd__or3b_1 _05397_ (.A(_00669_),
    .B(_01257_),
    .C_N(_00909_),
    .X(_01268_));
 sky130_fd_sc_hd__xnor2_1 _05398_ (.A(_00930_),
    .B(_01257_),
    .Y(net125));
 sky130_fd_sc_hd__and4_1 _05399_ (.A(net435),
    .B(net342),
    .C(net470),
    .D(net456),
    .X(_01289_));
 sky130_fd_sc_hd__a22oi_2 _05400_ (.A1(net342),
    .A2(net470),
    .B1(net456),
    .B2(net435),
    .Y(_01300_));
 sky130_fd_sc_hd__nand2_1 _05401_ (.A(net478),
    .B(net255),
    .Y(_01311_));
 sky130_fd_sc_hd__or3_1 _05402_ (.A(_01289_),
    .B(_01300_),
    .C(_01311_),
    .X(_01322_));
 sky130_fd_sc_hd__o21ai_1 _05403_ (.A1(_01289_),
    .A2(_01300_),
    .B1(_01311_),
    .Y(_01333_));
 sky130_fd_sc_hd__o21bai_1 _05404_ (.A1(_00962_),
    .A2(_00973_),
    .B1_N(_00951_),
    .Y(_01344_));
 sky130_fd_sc_hd__nand3_1 _05405_ (.A(_01322_),
    .B(_01333_),
    .C(_01344_),
    .Y(_01355_));
 sky130_fd_sc_hd__a21o_1 _05406_ (.A1(_01322_),
    .A2(_01333_),
    .B1(_01344_),
    .X(_01366_));
 sky130_fd_sc_hd__and4_1 _05407_ (.A(net485),
    .B(net493),
    .C(net235),
    .D(net227),
    .X(_01376_));
 sky130_fd_sc_hd__a22o_1 _05408_ (.A1(net485),
    .A2(net235),
    .B1(net227),
    .B2(net493),
    .X(_01387_));
 sky130_fd_sc_hd__and2b_1 _05409_ (.A_N(_01376_),
    .B(_01387_),
    .X(_01398_));
 sky130_fd_sc_hd__nand2_1 _05410_ (.A(net514),
    .B(net219),
    .Y(_01409_));
 sky130_fd_sc_hd__xnor2_1 _05411_ (.A(_01398_),
    .B(_01409_),
    .Y(_01420_));
 sky130_fd_sc_hd__nand3_1 _05412_ (.A(_01355_),
    .B(_01366_),
    .C(_01420_),
    .Y(_01431_));
 sky130_fd_sc_hd__a21o_1 _05413_ (.A1(_01355_),
    .A2(_01366_),
    .B1(_01420_),
    .X(_01442_));
 sky130_fd_sc_hd__a21bo_1 _05414_ (.A1(_01028_),
    .A2(_01082_),
    .B1_N(_01017_),
    .X(_01453_));
 sky130_fd_sc_hd__nand3_2 _05415_ (.A(_01431_),
    .B(_01442_),
    .C(_01453_),
    .Y(_01464_));
 sky130_fd_sc_hd__a21o_1 _05416_ (.A1(_01431_),
    .A2(_01442_),
    .B1(_01453_),
    .X(_01475_));
 sky130_fd_sc_hd__a31o_1 _05417_ (.A1(net599),
    .A2(net219),
    .A3(_01061_),
    .B1(_01039_),
    .X(_01486_));
 sky130_fd_sc_hd__and4_1 _05418_ (.A(net599),
    .B(net624),
    .C(net207),
    .D(net198),
    .X(_01497_));
 sky130_fd_sc_hd__a22oi_1 _05419_ (.A1(net599),
    .A2(net207),
    .B1(net198),
    .B2(net624),
    .Y(_01508_));
 sky130_fd_sc_hd__or2_1 _05420_ (.A(_01497_),
    .B(_01508_),
    .X(_01519_));
 sky130_fd_sc_hd__and2b_1 _05421_ (.A_N(_01519_),
    .B(_01486_),
    .X(_01529_));
 sky130_fd_sc_hd__xnor2_1 _05422_ (.A(_01486_),
    .B(_01519_),
    .Y(_01540_));
 sky130_fd_sc_hd__nand3_2 _05423_ (.A(_01464_),
    .B(_01475_),
    .C(_01540_),
    .Y(_01551_));
 sky130_fd_sc_hd__a21o_1 _05424_ (.A1(_01464_),
    .A2(_01475_),
    .B1(_01540_),
    .X(_01562_));
 sky130_fd_sc_hd__o211ai_4 _05425_ (.A1(_01126_),
    .A2(_01203_),
    .B1(_01551_),
    .C1(_01562_),
    .Y(_01573_));
 sky130_fd_sc_hd__a211o_1 _05426_ (.A1(_01551_),
    .A2(_01562_),
    .B1(_01126_),
    .C1(_01203_),
    .X(_01584_));
 sky130_fd_sc_hd__nand3_2 _05427_ (.A(_01181_),
    .B(_01573_),
    .C(_01584_),
    .Y(_01595_));
 sky130_fd_sc_hd__a21o_1 _05428_ (.A1(_01573_),
    .A2(_01584_),
    .B1(_01181_),
    .X(_01606_));
 sky130_fd_sc_hd__nand3_1 _05429_ (.A(_01246_),
    .B(_01595_),
    .C(_01606_),
    .Y(_01617_));
 sky130_fd_sc_hd__a21o_1 _05430_ (.A1(_01595_),
    .A2(_01606_),
    .B1(_01246_),
    .X(_01628_));
 sky130_fd_sc_hd__nand2_1 _05431_ (.A(_01617_),
    .B(_01628_),
    .Y(_01639_));
 sky130_fd_sc_hd__xor2_1 _05432_ (.A(_01268_),
    .B(_01639_),
    .X(net126));
 sky130_fd_sc_hd__or2_1 _05433_ (.A(_00669_),
    .B(_01257_),
    .X(_01660_));
 sky130_fd_sc_hd__nor3_2 _05434_ (.A(_00898_),
    .B(_01639_),
    .C(_01660_),
    .Y(_01671_));
 sky130_fd_sc_hd__and4bb_2 _05435_ (.A_N(_00778_),
    .B_N(_01660_),
    .C(_01628_),
    .D(_01617_),
    .X(_01682_));
 sky130_fd_sc_hd__nand2_1 _05436_ (.A(net255),
    .B(net470),
    .Y(_01693_));
 sky130_fd_sc_hd__and4_1 _05437_ (.A(net435),
    .B(net342),
    .C(net456),
    .D(net451),
    .X(_01703_));
 sky130_fd_sc_hd__a22oi_2 _05438_ (.A1(net342),
    .A2(net456),
    .B1(net451),
    .B2(net435),
    .Y(_01714_));
 sky130_fd_sc_hd__or3_1 _05439_ (.A(_01693_),
    .B(_01703_),
    .C(_01714_),
    .X(_01725_));
 sky130_fd_sc_hd__o21ai_1 _05440_ (.A1(_01703_),
    .A2(_01714_),
    .B1(_01693_),
    .Y(_01736_));
 sky130_fd_sc_hd__o21bai_1 _05441_ (.A1(_01300_),
    .A2(_01311_),
    .B1_N(_01289_),
    .Y(_01747_));
 sky130_fd_sc_hd__nand3_1 _05442_ (.A(_01725_),
    .B(_01736_),
    .C(_01747_),
    .Y(_01758_));
 sky130_fd_sc_hd__a21o_1 _05443_ (.A1(_01725_),
    .A2(_01736_),
    .B1(_01747_),
    .X(_01769_));
 sky130_fd_sc_hd__and4_1 _05444_ (.A(net478),
    .B(net485),
    .C(net236),
    .D(net227),
    .X(_01780_));
 sky130_fd_sc_hd__a22oi_1 _05445_ (.A1(net478),
    .A2(net236),
    .B1(net227),
    .B2(net485),
    .Y(_01791_));
 sky130_fd_sc_hd__nor2_1 _05446_ (.A(_01780_),
    .B(_01791_),
    .Y(_01802_));
 sky130_fd_sc_hd__nand2_1 _05447_ (.A(net493),
    .B(net219),
    .Y(_01813_));
 sky130_fd_sc_hd__xnor2_1 _05448_ (.A(_01802_),
    .B(_01813_),
    .Y(_01824_));
 sky130_fd_sc_hd__nand3_1 _05449_ (.A(_01758_),
    .B(_01769_),
    .C(_01824_),
    .Y(_01835_));
 sky130_fd_sc_hd__a21o_1 _05450_ (.A1(_01758_),
    .A2(_01769_),
    .B1(_01824_),
    .X(_01846_));
 sky130_fd_sc_hd__a21bo_1 _05451_ (.A1(_01366_),
    .A2(_01420_),
    .B1_N(_01355_),
    .X(_01857_));
 sky130_fd_sc_hd__and3_1 _05452_ (.A(_01835_),
    .B(_01846_),
    .C(_01857_),
    .X(_01867_));
 sky130_fd_sc_hd__a21oi_1 _05453_ (.A1(_01835_),
    .A2(_01846_),
    .B1(_01857_),
    .Y(_01878_));
 sky130_fd_sc_hd__a31o_1 _05454_ (.A1(net515),
    .A2(net219),
    .A3(_01387_),
    .B1(_01376_),
    .X(_01889_));
 sky130_fd_sc_hd__and4_1 _05455_ (.A(net515),
    .B(net599),
    .C(net207),
    .D(net198),
    .X(_01900_));
 sky130_fd_sc_hd__a22oi_1 _05456_ (.A1(net515),
    .A2(net207),
    .B1(net198),
    .B2(net599),
    .Y(_01911_));
 sky130_fd_sc_hd__nor2_1 _05457_ (.A(_01900_),
    .B(_01911_),
    .Y(_01922_));
 sky130_fd_sc_hd__nand2_1 _05458_ (.A(net624),
    .B(net196),
    .Y(_01933_));
 sky130_fd_sc_hd__xnor2_1 _05459_ (.A(_01922_),
    .B(_01933_),
    .Y(_01944_));
 sky130_fd_sc_hd__and2_1 _05460_ (.A(_01889_),
    .B(_01944_),
    .X(_01955_));
 sky130_fd_sc_hd__xor2_1 _05461_ (.A(_01889_),
    .B(_01944_),
    .X(_01966_));
 sky130_fd_sc_hd__and2_1 _05462_ (.A(_01497_),
    .B(_01966_),
    .X(_01977_));
 sky130_fd_sc_hd__xnor2_1 _05463_ (.A(_01497_),
    .B(_01966_),
    .Y(_01988_));
 sky130_fd_sc_hd__nor3_2 _05464_ (.A(_01867_),
    .B(_01878_),
    .C(_01988_),
    .Y(_01999_));
 sky130_fd_sc_hd__o21a_1 _05465_ (.A1(_01867_),
    .A2(_01878_),
    .B1(_01988_),
    .X(_02010_));
 sky130_fd_sc_hd__a211o_1 _05466_ (.A1(_01464_),
    .A2(_01551_),
    .B1(_01999_),
    .C1(_02010_),
    .X(_02021_));
 sky130_fd_sc_hd__o211ai_2 _05467_ (.A1(_01999_),
    .A2(_02010_),
    .B1(_01464_),
    .C1(_01551_),
    .Y(_02032_));
 sky130_fd_sc_hd__and3_1 _05468_ (.A(_01529_),
    .B(_02021_),
    .C(_02032_),
    .X(_02043_));
 sky130_fd_sc_hd__nand3_1 _05469_ (.A(_01529_),
    .B(_02021_),
    .C(_02032_),
    .Y(_02053_));
 sky130_fd_sc_hd__a21oi_1 _05470_ (.A1(_02021_),
    .A2(_02032_),
    .B1(_01529_),
    .Y(_02064_));
 sky130_fd_sc_hd__a211oi_2 _05471_ (.A1(_01573_),
    .A2(_01595_),
    .B1(_02043_),
    .C1(_02064_),
    .Y(_02075_));
 sky130_fd_sc_hd__o211a_1 _05472_ (.A1(_02043_),
    .A2(_02064_),
    .B1(_01573_),
    .C1(_01595_),
    .X(_02086_));
 sky130_fd_sc_hd__nor3_1 _05473_ (.A(_01617_),
    .B(_02075_),
    .C(_02086_),
    .Y(_02097_));
 sky130_fd_sc_hd__o21ai_1 _05474_ (.A1(_02075_),
    .A2(_02086_),
    .B1(_01617_),
    .Y(_02108_));
 sky130_fd_sc_hd__nand2b_1 _05475_ (.A_N(_02097_),
    .B(_02108_),
    .Y(_02119_));
 sky130_fd_sc_hd__xnor2_2 _05476_ (.A(_01682_),
    .B(_02119_),
    .Y(_02130_));
 sky130_fd_sc_hd__xor2_1 _05477_ (.A(_01671_),
    .B(_02130_),
    .X(net127));
 sky130_fd_sc_hd__o211a_1 _05478_ (.A1(_01955_),
    .A2(_01977_),
    .B1(net625),
    .C1(net187),
    .X(_02151_));
 sky130_fd_sc_hd__a211oi_1 _05479_ (.A1(net625),
    .A2(net187),
    .B1(_01955_),
    .C1(_01977_),
    .Y(_02162_));
 sky130_fd_sc_hd__nor2_1 _05480_ (.A(_02151_),
    .B(_02162_),
    .Y(_02173_));
 sky130_fd_sc_hd__o21ba_1 _05481_ (.A1(_01791_),
    .A2(_01813_),
    .B1_N(_01780_),
    .X(_02184_));
 sky130_fd_sc_hd__nand2_1 _05482_ (.A(net601),
    .B(net196),
    .Y(_02195_));
 sky130_fd_sc_hd__and4_1 _05483_ (.A(net493),
    .B(net515),
    .C(net207),
    .D(net198),
    .X(_02206_));
 sky130_fd_sc_hd__a22oi_1 _05484_ (.A1(net493),
    .A2(net207),
    .B1(net198),
    .B2(net515),
    .Y(_02216_));
 sky130_fd_sc_hd__nor2_1 _05485_ (.A(_02206_),
    .B(_02216_),
    .Y(_02227_));
 sky130_fd_sc_hd__xnor2_1 _05486_ (.A(_02195_),
    .B(_02227_),
    .Y(_02238_));
 sky130_fd_sc_hd__nand2b_1 _05487_ (.A_N(_02184_),
    .B(_02238_),
    .Y(_02249_));
 sky130_fd_sc_hd__xnor2_1 _05488_ (.A(_02184_),
    .B(_02238_),
    .Y(_02260_));
 sky130_fd_sc_hd__o21ba_1 _05489_ (.A1(_01911_),
    .A2(_01933_),
    .B1_N(_01900_),
    .X(_02271_));
 sky130_fd_sc_hd__nand2b_1 _05490_ (.A_N(_02271_),
    .B(_02260_),
    .Y(_02282_));
 sky130_fd_sc_hd__xnor2_1 _05491_ (.A(_02260_),
    .B(_02271_),
    .Y(_02293_));
 sky130_fd_sc_hd__and4_1 _05492_ (.A(net478),
    .B(net236),
    .C(net228),
    .D(net470),
    .X(_02304_));
 sky130_fd_sc_hd__a22oi_1 _05493_ (.A1(net478),
    .A2(net228),
    .B1(net470),
    .B2(net236),
    .Y(_02315_));
 sky130_fd_sc_hd__nor2_1 _05494_ (.A(_02304_),
    .B(_02315_),
    .Y(_02326_));
 sky130_fd_sc_hd__nand2_1 _05495_ (.A(net485),
    .B(net219),
    .Y(_02337_));
 sky130_fd_sc_hd__xnor2_1 _05496_ (.A(_02326_),
    .B(_02337_),
    .Y(_02348_));
 sky130_fd_sc_hd__nand2_1 _05497_ (.A(net255),
    .B(net456),
    .Y(_02359_));
 sky130_fd_sc_hd__and4_1 _05498_ (.A(net435),
    .B(net342),
    .C(net451),
    .D(net445),
    .X(_02370_));
 sky130_fd_sc_hd__a22oi_2 _05499_ (.A1(net342),
    .A2(net451),
    .B1(net445),
    .B2(net435),
    .Y(_02380_));
 sky130_fd_sc_hd__or3_1 _05500_ (.A(_02359_),
    .B(_02370_),
    .C(_02380_),
    .X(_02391_));
 sky130_fd_sc_hd__o21ai_1 _05501_ (.A1(_02370_),
    .A2(_02380_),
    .B1(_02359_),
    .Y(_02402_));
 sky130_fd_sc_hd__o21bai_1 _05502_ (.A1(_01693_),
    .A2(_01714_),
    .B1_N(_01703_),
    .Y(_02413_));
 sky130_fd_sc_hd__nand3_1 _05503_ (.A(_02391_),
    .B(_02402_),
    .C(_02413_),
    .Y(_02424_));
 sky130_fd_sc_hd__a21o_1 _05504_ (.A1(_02391_),
    .A2(_02402_),
    .B1(_02413_),
    .X(_02435_));
 sky130_fd_sc_hd__nand3_1 _05505_ (.A(_02348_),
    .B(_02424_),
    .C(_02435_),
    .Y(_02446_));
 sky130_fd_sc_hd__a21o_1 _05506_ (.A1(_02424_),
    .A2(_02435_),
    .B1(_02348_),
    .X(_02457_));
 sky130_fd_sc_hd__a21bo_1 _05507_ (.A1(_01769_),
    .A2(_01824_),
    .B1_N(_01758_),
    .X(_02468_));
 sky130_fd_sc_hd__nand3_2 _05508_ (.A(_02446_),
    .B(_02457_),
    .C(_02468_),
    .Y(_02479_));
 sky130_fd_sc_hd__a21o_1 _05509_ (.A1(_02446_),
    .A2(_02457_),
    .B1(_02468_),
    .X(_02490_));
 sky130_fd_sc_hd__nand3_2 _05510_ (.A(_02293_),
    .B(_02479_),
    .C(_02490_),
    .Y(_02501_));
 sky130_fd_sc_hd__a21o_1 _05511_ (.A1(_02479_),
    .A2(_02490_),
    .B1(_02293_),
    .X(_02512_));
 sky130_fd_sc_hd__o211a_1 _05512_ (.A1(_01867_),
    .A2(_01999_),
    .B1(_02501_),
    .C1(_02512_),
    .X(_02523_));
 sky130_fd_sc_hd__o211ai_1 _05513_ (.A1(_01867_),
    .A2(_01999_),
    .B1(_02501_),
    .C1(_02512_),
    .Y(_02534_));
 sky130_fd_sc_hd__a211o_1 _05514_ (.A1(_02501_),
    .A2(_02512_),
    .B1(_01867_),
    .C1(_01999_),
    .X(_02544_));
 sky130_fd_sc_hd__and3_1 _05515_ (.A(_02173_),
    .B(_02534_),
    .C(_02544_),
    .X(_02555_));
 sky130_fd_sc_hd__a21oi_1 _05516_ (.A1(_02534_),
    .A2(_02544_),
    .B1(_02173_),
    .Y(_02566_));
 sky130_fd_sc_hd__a211o_1 _05517_ (.A1(_02021_),
    .A2(_02053_),
    .B1(_02555_),
    .C1(_02566_),
    .X(_02577_));
 sky130_fd_sc_hd__o211ai_1 _05518_ (.A1(_02555_),
    .A2(_02566_),
    .B1(_02021_),
    .C1(_02053_),
    .Y(_02588_));
 sky130_fd_sc_hd__and3_1 _05519_ (.A(_02075_),
    .B(_02577_),
    .C(_02588_),
    .X(_02599_));
 sky130_fd_sc_hd__inv_2 _05520_ (.A(_02599_),
    .Y(_02610_));
 sky130_fd_sc_hd__a21o_1 _05521_ (.A1(_02577_),
    .A2(_02588_),
    .B1(_02075_),
    .X(_02621_));
 sky130_fd_sc_hd__and2b_1 _05522_ (.A_N(_02599_),
    .B(_02621_),
    .X(_02632_));
 sky130_fd_sc_hd__nand4b_1 _05523_ (.A_N(net142),
    .B(_02108_),
    .C(_02632_),
    .D(_01682_),
    .Y(_02643_));
 sky130_fd_sc_hd__o21ba_1 _05524_ (.A1(_02195_),
    .A2(_02216_),
    .B1_N(_02206_),
    .X(_02654_));
 sky130_fd_sc_hd__o21ba_1 _05525_ (.A1(_02315_),
    .A2(_02337_),
    .B1_N(_02304_),
    .X(_02665_));
 sky130_fd_sc_hd__and4_1 _05526_ (.A(net486),
    .B(net493),
    .C(net207),
    .D(net198),
    .X(_02676_));
 sky130_fd_sc_hd__a22oi_1 _05527_ (.A1(net486),
    .A2(net207),
    .B1(net198),
    .B2(net493),
    .Y(_02687_));
 sky130_fd_sc_hd__nor2_1 _05528_ (.A(_02676_),
    .B(_02687_),
    .Y(_02697_));
 sky130_fd_sc_hd__nand2_1 _05529_ (.A(net515),
    .B(net196),
    .Y(_02708_));
 sky130_fd_sc_hd__xnor2_1 _05530_ (.A(_02697_),
    .B(_02708_),
    .Y(_02719_));
 sky130_fd_sc_hd__nand2b_1 _05531_ (.A_N(_02665_),
    .B(_02719_),
    .Y(_02730_));
 sky130_fd_sc_hd__xnor2_1 _05532_ (.A(_02665_),
    .B(_02719_),
    .Y(_02741_));
 sky130_fd_sc_hd__nand2b_1 _05533_ (.A_N(_02654_),
    .B(_02741_),
    .Y(_02752_));
 sky130_fd_sc_hd__xnor2_1 _05534_ (.A(_02654_),
    .B(_02741_),
    .Y(_02763_));
 sky130_fd_sc_hd__and4_1 _05535_ (.A(net236),
    .B(net228),
    .C(net470),
    .D(net456),
    .X(_02774_));
 sky130_fd_sc_hd__a22oi_1 _05536_ (.A1(net228),
    .A2(net470),
    .B1(net456),
    .B2(net236),
    .Y(_02785_));
 sky130_fd_sc_hd__nor2_1 _05537_ (.A(_02774_),
    .B(_02785_),
    .Y(_02796_));
 sky130_fd_sc_hd__nand2_1 _05538_ (.A(net478),
    .B(net219),
    .Y(_02807_));
 sky130_fd_sc_hd__xnor2_1 _05539_ (.A(_02796_),
    .B(_02807_),
    .Y(_02818_));
 sky130_fd_sc_hd__nand2_1 _05540_ (.A(net255),
    .B(net451),
    .Y(_02829_));
 sky130_fd_sc_hd__and4_1 _05541_ (.A(net435),
    .B(net342),
    .C(net546),
    .D(net445),
    .X(_02840_));
 sky130_fd_sc_hd__a22oi_2 _05542_ (.A1(net441),
    .A2(net546),
    .B1(net445),
    .B2(net44),
    .Y(_02850_));
 sky130_fd_sc_hd__or3_1 _05543_ (.A(_02829_),
    .B(_02840_),
    .C(_02850_),
    .X(_02861_));
 sky130_fd_sc_hd__o21ai_1 _05544_ (.A1(_02840_),
    .A2(_02850_),
    .B1(_02829_),
    .Y(_02872_));
 sky130_fd_sc_hd__o21bai_1 _05545_ (.A1(_02359_),
    .A2(_02380_),
    .B1_N(_02370_),
    .Y(_02883_));
 sky130_fd_sc_hd__nand3_1 _05546_ (.A(_02861_),
    .B(_02872_),
    .C(_02883_),
    .Y(_02894_));
 sky130_fd_sc_hd__a21o_1 _05547_ (.A1(_02861_),
    .A2(_02872_),
    .B1(_02883_),
    .X(_02905_));
 sky130_fd_sc_hd__nand3_1 _05548_ (.A(_02818_),
    .B(_02894_),
    .C(_02905_),
    .Y(_02916_));
 sky130_fd_sc_hd__a21o_1 _05549_ (.A1(_02894_),
    .A2(_02905_),
    .B1(_02818_),
    .X(_02927_));
 sky130_fd_sc_hd__a21bo_1 _05550_ (.A1(_02348_),
    .A2(_02435_),
    .B1_N(_02424_),
    .X(_02938_));
 sky130_fd_sc_hd__nand3_2 _05551_ (.A(_02916_),
    .B(_02927_),
    .C(_02938_),
    .Y(_02949_));
 sky130_fd_sc_hd__a21o_1 _05552_ (.A1(_02916_),
    .A2(_02927_),
    .B1(_02938_),
    .X(_02960_));
 sky130_fd_sc_hd__and3_1 _05553_ (.A(_02763_),
    .B(_02949_),
    .C(_02960_),
    .X(_02971_));
 sky130_fd_sc_hd__nand3_1 _05554_ (.A(_02763_),
    .B(_02949_),
    .C(_02960_),
    .Y(_02982_));
 sky130_fd_sc_hd__a21oi_1 _05555_ (.A1(_02949_),
    .A2(_02960_),
    .B1(_02763_),
    .Y(_02993_));
 sky130_fd_sc_hd__a211o_1 _05556_ (.A1(_02479_),
    .A2(_02501_),
    .B1(_02971_),
    .C1(_02993_),
    .X(_03003_));
 sky130_fd_sc_hd__o211ai_2 _05557_ (.A1(_02971_),
    .A2(_02993_),
    .B1(_02479_),
    .C1(_02501_),
    .Y(_03014_));
 sky130_fd_sc_hd__a22oi_1 _05558_ (.A1(net601),
    .A2(net187),
    .B1(net430),
    .B2(net625),
    .Y(_03025_));
 sky130_fd_sc_hd__and4_1 _05559_ (.A(net601),
    .B(net625),
    .C(net187),
    .D(net430),
    .X(_03036_));
 sky130_fd_sc_hd__or2_1 _05560_ (.A(_03025_),
    .B(_03036_),
    .X(_03047_));
 sky130_fd_sc_hd__a21oi_1 _05561_ (.A1(_02249_),
    .A2(_02282_),
    .B1(_03047_),
    .Y(_03058_));
 sky130_fd_sc_hd__and3_1 _05562_ (.A(_02249_),
    .B(_02282_),
    .C(_03047_),
    .X(_03069_));
 sky130_fd_sc_hd__nor2_1 _05563_ (.A(_03058_),
    .B(_03069_),
    .Y(_03080_));
 sky130_fd_sc_hd__nand3_2 _05564_ (.A(_03003_),
    .B(_03014_),
    .C(_03080_),
    .Y(_03091_));
 sky130_fd_sc_hd__a21o_1 _05565_ (.A1(_03003_),
    .A2(_03014_),
    .B1(_03080_),
    .X(_03102_));
 sky130_fd_sc_hd__o211ai_1 _05566_ (.A1(_02523_),
    .A2(_02555_),
    .B1(_03091_),
    .C1(_03102_),
    .Y(_03113_));
 sky130_fd_sc_hd__a211o_1 _05567_ (.A1(_03091_),
    .A2(_03102_),
    .B1(_02523_),
    .C1(_02555_),
    .X(_03124_));
 sky130_fd_sc_hd__and3_1 _05568_ (.A(_02151_),
    .B(_03113_),
    .C(_03124_),
    .X(_03134_));
 sky130_fd_sc_hd__a21oi_1 _05569_ (.A1(_03113_),
    .A2(_03124_),
    .B1(_02151_),
    .Y(_03145_));
 sky130_fd_sc_hd__or3_2 _05570_ (.A(_02577_),
    .B(_03134_),
    .C(_03145_),
    .X(_03156_));
 sky130_fd_sc_hd__o21ai_2 _05571_ (.A1(_03134_),
    .A2(_03145_),
    .B1(_02577_),
    .Y(_03167_));
 sky130_fd_sc_hd__a21oi_1 _05572_ (.A1(net142),
    .A2(_02621_),
    .B1(_02599_),
    .Y(_03178_));
 sky130_fd_sc_hd__nand3_1 _05573_ (.A(_03156_),
    .B(_03167_),
    .C(_03178_),
    .Y(_03189_));
 sky130_fd_sc_hd__a21o_1 _05574_ (.A1(_03156_),
    .A2(_03167_),
    .B1(_03178_),
    .X(_03200_));
 sky130_fd_sc_hd__a21oi_1 _05575_ (.A1(_03189_),
    .A2(_03200_),
    .B1(_02643_),
    .Y(_03211_));
 sky130_fd_sc_hd__and3_1 _05576_ (.A(_02643_),
    .B(_03189_),
    .C(_03200_),
    .X(_03222_));
 sky130_fd_sc_hd__nor2_1 _05577_ (.A(_03211_),
    .B(_03222_),
    .Y(_03233_));
 sky130_fd_sc_hd__a21oi_1 _05578_ (.A1(_01682_),
    .A2(_02108_),
    .B1(_02097_),
    .Y(_03244_));
 sky130_fd_sc_hd__xnor2_1 _05579_ (.A(_02632_),
    .B(_03244_),
    .Y(_03255_));
 sky130_fd_sc_hd__and3_1 _05580_ (.A(_01671_),
    .B(_02130_),
    .C(_03255_),
    .X(_03266_));
 sky130_fd_sc_hd__nand3_1 _05581_ (.A(_01671_),
    .B(_02130_),
    .C(_03255_),
    .Y(_03276_));
 sky130_fd_sc_hd__xnor2_1 _05582_ (.A(_03233_),
    .B(_03276_),
    .Y(net66));
 sky130_fd_sc_hd__and4_1 _05583_ (.A(net142),
    .B(_02632_),
    .C(_03156_),
    .D(_03167_),
    .X(_03297_));
 sky130_fd_sc_hd__and4_1 _05584_ (.A(net515),
    .B(net600),
    .C(net187),
    .D(net430),
    .X(_03308_));
 sky130_fd_sc_hd__a22oi_1 _05585_ (.A1(net515),
    .A2(net187),
    .B1(net430),
    .B2(net600),
    .Y(_03319_));
 sky130_fd_sc_hd__nor2_1 _05586_ (.A(_03308_),
    .B(_03319_),
    .Y(_03330_));
 sky130_fd_sc_hd__nand2_1 _05587_ (.A(net625),
    .B(net423),
    .Y(_03341_));
 sky130_fd_sc_hd__xnor2_1 _05588_ (.A(_03330_),
    .B(_03341_),
    .Y(_03352_));
 sky130_fd_sc_hd__and2_1 _05589_ (.A(_03036_),
    .B(_03352_),
    .X(_03363_));
 sky130_fd_sc_hd__nor2_1 _05590_ (.A(_03036_),
    .B(_03352_),
    .Y(_03374_));
 sky130_fd_sc_hd__or2_1 _05591_ (.A(_03363_),
    .B(_03374_),
    .X(_03385_));
 sky130_fd_sc_hd__a21oi_1 _05592_ (.A1(_02730_),
    .A2(_02752_),
    .B1(_03385_),
    .Y(_03395_));
 sky130_fd_sc_hd__and3_1 _05593_ (.A(_02730_),
    .B(_02752_),
    .C(_03385_),
    .X(_03406_));
 sky130_fd_sc_hd__nor2_1 _05594_ (.A(_03395_),
    .B(_03406_),
    .Y(_03417_));
 sky130_fd_sc_hd__o21ba_1 _05595_ (.A1(_02687_),
    .A2(_02708_),
    .B1_N(_02676_),
    .X(_03428_));
 sky130_fd_sc_hd__o21ba_1 _05596_ (.A1(_02785_),
    .A2(_02807_),
    .B1_N(_02774_),
    .X(_03439_));
 sky130_fd_sc_hd__and4_1 _05597_ (.A(net479),
    .B(net486),
    .C(net208),
    .D(net198),
    .X(_03450_));
 sky130_fd_sc_hd__a22oi_1 _05598_ (.A1(net479),
    .A2(net208),
    .B1(net198),
    .B2(net486),
    .Y(_03461_));
 sky130_fd_sc_hd__nor2_1 _05599_ (.A(_03450_),
    .B(_03461_),
    .Y(_03472_));
 sky130_fd_sc_hd__nand2_1 _05600_ (.A(net493),
    .B(net196),
    .Y(_03483_));
 sky130_fd_sc_hd__xnor2_1 _05601_ (.A(_03472_),
    .B(_03483_),
    .Y(_03494_));
 sky130_fd_sc_hd__nand2b_1 _05602_ (.A_N(_03439_),
    .B(_03494_),
    .Y(_03505_));
 sky130_fd_sc_hd__xnor2_1 _05603_ (.A(_03439_),
    .B(_03494_),
    .Y(_03515_));
 sky130_fd_sc_hd__nand2b_1 _05604_ (.A_N(_03428_),
    .B(_03515_),
    .Y(_03526_));
 sky130_fd_sc_hd__xnor2_1 _05605_ (.A(_03428_),
    .B(_03515_),
    .Y(_03537_));
 sky130_fd_sc_hd__nand2_1 _05606_ (.A(net219),
    .B(net470),
    .Y(_03548_));
 sky130_fd_sc_hd__and4_1 _05607_ (.A(net236),
    .B(net228),
    .C(net456),
    .D(net451),
    .X(_03559_));
 sky130_fd_sc_hd__a22oi_1 _05608_ (.A1(net228),
    .A2(net456),
    .B1(net451),
    .B2(net236),
    .Y(_03570_));
 sky130_fd_sc_hd__nor2_1 _05609_ (.A(_03559_),
    .B(_03570_),
    .Y(_03581_));
 sky130_fd_sc_hd__xnor2_1 _05610_ (.A(_03548_),
    .B(_03581_),
    .Y(_03592_));
 sky130_fd_sc_hd__nand2_1 _05611_ (.A(net258),
    .B(net445),
    .Y(_03603_));
 sky130_fd_sc_hd__and4_1 _05612_ (.A(net440),
    .B(net347),
    .C(net546),
    .D(net465),
    .X(_03614_));
 sky130_fd_sc_hd__a22oi_2 _05613_ (.A1(net347),
    .A2(net546),
    .B1(net465),
    .B2(net440),
    .Y(_03624_));
 sky130_fd_sc_hd__or3_1 _05614_ (.A(_03603_),
    .B(_03614_),
    .C(_03624_),
    .X(_03635_));
 sky130_fd_sc_hd__o21ai_1 _05615_ (.A1(_03614_),
    .A2(_03624_),
    .B1(_03603_),
    .Y(_03646_));
 sky130_fd_sc_hd__o21bai_1 _05616_ (.A1(_02829_),
    .A2(_02850_),
    .B1_N(_02840_),
    .Y(_03657_));
 sky130_fd_sc_hd__nand3_1 _05617_ (.A(_03635_),
    .B(_03646_),
    .C(_03657_),
    .Y(_03668_));
 sky130_fd_sc_hd__a21o_1 _05618_ (.A1(_03635_),
    .A2(_03646_),
    .B1(_03657_),
    .X(_03679_));
 sky130_fd_sc_hd__nand3_1 _05619_ (.A(_03592_),
    .B(_03668_),
    .C(_03679_),
    .Y(_03690_));
 sky130_fd_sc_hd__a21o_1 _05620_ (.A1(_03668_),
    .A2(_03679_),
    .B1(_03592_),
    .X(_03701_));
 sky130_fd_sc_hd__a21bo_1 _05621_ (.A1(_02818_),
    .A2(_02905_),
    .B1_N(_02894_),
    .X(_03712_));
 sky130_fd_sc_hd__nand3_1 _05622_ (.A(_03690_),
    .B(_03701_),
    .C(_03712_),
    .Y(_03723_));
 sky130_fd_sc_hd__inv_2 _05623_ (.A(_03723_),
    .Y(_03734_));
 sky130_fd_sc_hd__a21o_1 _05624_ (.A1(_03690_),
    .A2(_03701_),
    .B1(_03712_),
    .X(_03744_));
 sky130_fd_sc_hd__and3_1 _05625_ (.A(_03537_),
    .B(_03723_),
    .C(_03744_),
    .X(_03755_));
 sky130_fd_sc_hd__a21oi_1 _05626_ (.A1(_03723_),
    .A2(_03744_),
    .B1(_03537_),
    .Y(_03766_));
 sky130_fd_sc_hd__a211o_1 _05627_ (.A1(_02949_),
    .A2(_02982_),
    .B1(_03755_),
    .C1(_03766_),
    .X(_03777_));
 sky130_fd_sc_hd__o211ai_2 _05628_ (.A1(_03755_),
    .A2(_03766_),
    .B1(_02949_),
    .C1(_02982_),
    .Y(_03788_));
 sky130_fd_sc_hd__and3_1 _05629_ (.A(_03417_),
    .B(_03777_),
    .C(_03788_),
    .X(_03799_));
 sky130_fd_sc_hd__a21oi_1 _05630_ (.A1(_03777_),
    .A2(_03788_),
    .B1(_03417_),
    .Y(_03810_));
 sky130_fd_sc_hd__a211o_2 _05631_ (.A1(_03003_),
    .A2(_03091_),
    .B1(_03799_),
    .C1(_03810_),
    .X(_03821_));
 sky130_fd_sc_hd__o211ai_2 _05632_ (.A1(_03799_),
    .A2(_03810_),
    .B1(_03003_),
    .C1(_03091_),
    .Y(_03832_));
 sky130_fd_sc_hd__nand3_2 _05633_ (.A(_03058_),
    .B(_03821_),
    .C(_03832_),
    .Y(_03843_));
 sky130_fd_sc_hd__a21o_1 _05634_ (.A1(_03821_),
    .A2(_03832_),
    .B1(_03058_),
    .X(_03853_));
 sky130_fd_sc_hd__and2_1 _05635_ (.A(_03843_),
    .B(_03853_),
    .X(_03864_));
 sky130_fd_sc_hd__a21bo_1 _05636_ (.A1(_02151_),
    .A2(_03124_),
    .B1_N(_03113_),
    .X(_03875_));
 sky130_fd_sc_hd__nand2_1 _05637_ (.A(_03864_),
    .B(_03875_),
    .Y(_03886_));
 sky130_fd_sc_hd__xnor2_1 _05638_ (.A(_03864_),
    .B(_03875_),
    .Y(_03897_));
 sky130_fd_sc_hd__a21bo_1 _05639_ (.A1(_02599_),
    .A2(_03167_),
    .B1_N(_03156_),
    .X(_03908_));
 sky130_fd_sc_hd__nor2_1 _05640_ (.A(_03156_),
    .B(_03897_),
    .Y(_03919_));
 sky130_fd_sc_hd__and4bb_1 _05641_ (.A_N(_02610_),
    .B_N(_03897_),
    .C(_03167_),
    .D(_03156_),
    .X(_03930_));
 sky130_fd_sc_hd__xnor2_1 _05642_ (.A(_03897_),
    .B(_03908_),
    .Y(_03941_));
 sky130_fd_sc_hd__and2_1 _05643_ (.A(_03297_),
    .B(_03941_),
    .X(_03951_));
 sky130_fd_sc_hd__xor2_1 _05644_ (.A(_03297_),
    .B(_03941_),
    .X(_03962_));
 sky130_fd_sc_hd__o21bai_1 _05645_ (.A1(_03222_),
    .A2(_03276_),
    .B1_N(_03211_),
    .Y(_03973_));
 sky130_fd_sc_hd__xor2_1 _05646_ (.A(_03962_),
    .B(_03973_),
    .X(net67));
 sky130_fd_sc_hd__nand2_1 _05647_ (.A(_03505_),
    .B(_03526_),
    .Y(_03994_));
 sky130_fd_sc_hd__and4_1 _05648_ (.A(net493),
    .B(net516),
    .C(net187),
    .D(net430),
    .X(_04005_));
 sky130_fd_sc_hd__a22oi_1 _05649_ (.A1(net494),
    .A2(net187),
    .B1(net430),
    .B2(net516),
    .Y(_04016_));
 sky130_fd_sc_hd__nor2_1 _05650_ (.A(_04005_),
    .B(_04016_),
    .Y(_04027_));
 sky130_fd_sc_hd__nand2_1 _05651_ (.A(net600),
    .B(net423),
    .Y(_04038_));
 sky130_fd_sc_hd__xnor2_1 _05652_ (.A(_04027_),
    .B(_04038_),
    .Y(_04048_));
 sky130_fd_sc_hd__o21ba_1 _05653_ (.A1(_03319_),
    .A2(_03341_),
    .B1_N(_03308_),
    .X(_04059_));
 sky130_fd_sc_hd__nand2b_1 _05654_ (.A_N(_04059_),
    .B(_04048_),
    .Y(_04070_));
 sky130_fd_sc_hd__xnor2_1 _05655_ (.A(_04048_),
    .B(_04059_),
    .Y(_04081_));
 sky130_fd_sc_hd__nand3_2 _05656_ (.A(net625),
    .B(net419),
    .C(_04081_),
    .Y(_04092_));
 sky130_fd_sc_hd__a21o_1 _05657_ (.A1(net625),
    .A2(net419),
    .B1(_04081_),
    .X(_04103_));
 sky130_fd_sc_hd__nand2_1 _05658_ (.A(_04092_),
    .B(_04103_),
    .Y(_04114_));
 sky130_fd_sc_hd__xnor2_1 _05659_ (.A(_03994_),
    .B(_04114_),
    .Y(_04125_));
 sky130_fd_sc_hd__xnor2_1 _05660_ (.A(_03363_),
    .B(_04125_),
    .Y(_04136_));
 sky130_fd_sc_hd__o21ba_1 _05661_ (.A1(_03461_),
    .A2(_03483_),
    .B1_N(_03450_),
    .X(_04146_));
 sky130_fd_sc_hd__o21ba_1 _05662_ (.A1(_03548_),
    .A2(_03570_),
    .B1_N(_03559_),
    .X(_04157_));
 sky130_fd_sc_hd__and4_1 _05663_ (.A(net479),
    .B(net471),
    .C(net208),
    .D(net199),
    .X(_04168_));
 sky130_fd_sc_hd__a22oi_1 _05664_ (.A1(net471),
    .A2(net208),
    .B1(net199),
    .B2(net479),
    .Y(_04179_));
 sky130_fd_sc_hd__nor2_1 _05665_ (.A(_04168_),
    .B(_04179_),
    .Y(_04190_));
 sky130_fd_sc_hd__nand2_1 _05666_ (.A(net486),
    .B(net196),
    .Y(_04201_));
 sky130_fd_sc_hd__xnor2_1 _05667_ (.A(_04190_),
    .B(_04201_),
    .Y(_04212_));
 sky130_fd_sc_hd__and2b_1 _05668_ (.A_N(_04157_),
    .B(_04212_),
    .X(_04223_));
 sky130_fd_sc_hd__xnor2_1 _05669_ (.A(_04157_),
    .B(_04212_),
    .Y(_04233_));
 sky130_fd_sc_hd__and2b_1 _05670_ (.A_N(_04146_),
    .B(_04233_),
    .X(_04244_));
 sky130_fd_sc_hd__xnor2_1 _05671_ (.A(_04146_),
    .B(_04233_),
    .Y(_04255_));
 sky130_fd_sc_hd__nand2_1 _05672_ (.A(net219),
    .B(net456),
    .Y(_04266_));
 sky130_fd_sc_hd__and4_1 _05673_ (.A(net242),
    .B(net234),
    .C(net451),
    .D(net445),
    .X(_04277_));
 sky130_fd_sc_hd__a22oi_1 _05674_ (.A1(net228),
    .A2(net451),
    .B1(net445),
    .B2(net242),
    .Y(_04288_));
 sky130_fd_sc_hd__nor2_1 _05675_ (.A(_04277_),
    .B(_04288_),
    .Y(_04299_));
 sky130_fd_sc_hd__xnor2_1 _05676_ (.A(_04266_),
    .B(_04299_),
    .Y(_04310_));
 sky130_fd_sc_hd__nand2_1 _05677_ (.A(net256),
    .B(net546),
    .Y(_04320_));
 sky130_fd_sc_hd__and4_1 _05678_ (.A(net440),
    .B(net347),
    .C(net465),
    .D(net384),
    .X(_04331_));
 sky130_fd_sc_hd__a22oi_2 _05679_ (.A1(net347),
    .A2(net465),
    .B1(net384),
    .B2(net440),
    .Y(_04342_));
 sky130_fd_sc_hd__or3_1 _05680_ (.A(_04320_),
    .B(_04331_),
    .C(_04342_),
    .X(_04353_));
 sky130_fd_sc_hd__o21ai_1 _05681_ (.A1(_04331_),
    .A2(_04342_),
    .B1(_04320_),
    .Y(_04364_));
 sky130_fd_sc_hd__o21bai_1 _05682_ (.A1(_03603_),
    .A2(_03624_),
    .B1_N(_03614_),
    .Y(_04375_));
 sky130_fd_sc_hd__nand3_1 _05683_ (.A(_04353_),
    .B(_04364_),
    .C(_04375_),
    .Y(_04385_));
 sky130_fd_sc_hd__a21o_1 _05684_ (.A1(_04353_),
    .A2(_04364_),
    .B1(_04375_),
    .X(_04396_));
 sky130_fd_sc_hd__nand3_1 _05685_ (.A(_04310_),
    .B(_04385_),
    .C(_04396_),
    .Y(_04407_));
 sky130_fd_sc_hd__a21o_1 _05686_ (.A1(_04385_),
    .A2(_04396_),
    .B1(_04310_),
    .X(_04418_));
 sky130_fd_sc_hd__a21bo_1 _05687_ (.A1(_03592_),
    .A2(_03679_),
    .B1_N(_03668_),
    .X(_04429_));
 sky130_fd_sc_hd__nand3_2 _05688_ (.A(_04407_),
    .B(_04418_),
    .C(_04429_),
    .Y(_04440_));
 sky130_fd_sc_hd__a21o_1 _05689_ (.A1(_04407_),
    .A2(_04418_),
    .B1(_04429_),
    .X(_04451_));
 sky130_fd_sc_hd__nand3_1 _05690_ (.A(_04255_),
    .B(_04440_),
    .C(_04451_),
    .Y(_04461_));
 sky130_fd_sc_hd__a21o_1 _05691_ (.A1(_04440_),
    .A2(_04451_),
    .B1(_04255_),
    .X(_04472_));
 sky130_fd_sc_hd__o211a_1 _05692_ (.A1(_03734_),
    .A2(_03755_),
    .B1(_04461_),
    .C1(_04472_),
    .X(_04483_));
 sky130_fd_sc_hd__a211oi_1 _05693_ (.A1(_04461_),
    .A2(_04472_),
    .B1(_03734_),
    .C1(_03755_),
    .Y(_04494_));
 sky130_fd_sc_hd__nor2_1 _05694_ (.A(_04483_),
    .B(_04494_),
    .Y(_04505_));
 sky130_fd_sc_hd__xnor2_1 _05695_ (.A(_04136_),
    .B(_04505_),
    .Y(_04516_));
 sky130_fd_sc_hd__a21bo_1 _05696_ (.A1(_03417_),
    .A2(_03788_),
    .B1_N(_03777_),
    .X(_04526_));
 sky130_fd_sc_hd__and2_1 _05697_ (.A(_04516_),
    .B(_04526_),
    .X(_04537_));
 sky130_fd_sc_hd__xor2_1 _05698_ (.A(_04516_),
    .B(_04526_),
    .X(_04548_));
 sky130_fd_sc_hd__and2_1 _05699_ (.A(_03395_),
    .B(_04548_),
    .X(_04559_));
 sky130_fd_sc_hd__nor2_1 _05700_ (.A(_03395_),
    .B(_04548_),
    .Y(_04570_));
 sky130_fd_sc_hd__a211oi_4 _05701_ (.A1(_03821_),
    .A2(_03843_),
    .B1(_04559_),
    .C1(_04570_),
    .Y(_04581_));
 sky130_fd_sc_hd__o211a_1 _05702_ (.A1(_04559_),
    .A2(_04570_),
    .B1(_03821_),
    .C1(_03843_),
    .X(_04591_));
 sky130_fd_sc_hd__or3_1 _05703_ (.A(_03886_),
    .B(_04581_),
    .C(_04591_),
    .X(_04602_));
 sky130_fd_sc_hd__o21ai_1 _05704_ (.A1(_04581_),
    .A2(_04591_),
    .B1(_03886_),
    .Y(_04613_));
 sky130_fd_sc_hd__nand3_2 _05705_ (.A(_03919_),
    .B(_04602_),
    .C(_04613_),
    .Y(_04624_));
 sky130_fd_sc_hd__a21o_1 _05706_ (.A1(_04602_),
    .A2(_04613_),
    .B1(_03919_),
    .X(_04635_));
 sky130_fd_sc_hd__and3_1 _05707_ (.A(_03930_),
    .B(_04624_),
    .C(_04635_),
    .X(_04645_));
 sky130_fd_sc_hd__a21o_1 _05708_ (.A1(_04624_),
    .A2(_04635_),
    .B1(_03930_),
    .X(_04656_));
 sky130_fd_sc_hd__nand2b_1 _05709_ (.A_N(_04645_),
    .B(_04656_),
    .Y(_04667_));
 sky130_fd_sc_hd__a21o_1 _05710_ (.A1(_03962_),
    .A2(_03973_),
    .B1(_03951_),
    .X(_04678_));
 sky130_fd_sc_hd__xnor2_1 _05711_ (.A(_04667_),
    .B(_04678_),
    .Y(net68));
 sky130_fd_sc_hd__a21oi_1 _05712_ (.A1(_04656_),
    .A2(_04678_),
    .B1(_04645_),
    .Y(_04698_));
 sky130_fd_sc_hd__a32oi_2 _05713_ (.A1(_03994_),
    .A2(_04092_),
    .A3(_04103_),
    .B1(_04125_),
    .B2(_03363_),
    .Y(_04709_));
 sky130_fd_sc_hd__a22oi_1 _05714_ (.A1(net600),
    .A2(net419),
    .B1(net411),
    .B2(net625),
    .Y(_04720_));
 sky130_fd_sc_hd__and4_1 _05715_ (.A(net600),
    .B(net625),
    .C(net419),
    .D(net411),
    .X(_04730_));
 sky130_fd_sc_hd__or2_1 _05716_ (.A(_04720_),
    .B(_04730_),
    .X(_04741_));
 sky130_fd_sc_hd__and4_1 _05717_ (.A(net487),
    .B(net495),
    .C(net187),
    .D(net430),
    .X(_04752_));
 sky130_fd_sc_hd__a22oi_1 _05718_ (.A1(net487),
    .A2(net187),
    .B1(net430),
    .B2(net495),
    .Y(_04763_));
 sky130_fd_sc_hd__nor2_1 _05719_ (.A(_04752_),
    .B(_04763_),
    .Y(_04773_));
 sky130_fd_sc_hd__nand2_1 _05720_ (.A(net516),
    .B(net423),
    .Y(_04784_));
 sky130_fd_sc_hd__xnor2_1 _05721_ (.A(_04773_),
    .B(_04784_),
    .Y(_04795_));
 sky130_fd_sc_hd__o21ba_1 _05722_ (.A1(_04016_),
    .A2(_04038_),
    .B1_N(_04005_),
    .X(_04805_));
 sky130_fd_sc_hd__nand2b_1 _05723_ (.A_N(_04805_),
    .B(_04795_),
    .Y(_04816_));
 sky130_fd_sc_hd__xnor2_1 _05724_ (.A(_04795_),
    .B(_04805_),
    .Y(_04826_));
 sky130_fd_sc_hd__nand2b_1 _05725_ (.A_N(_04741_),
    .B(_04826_),
    .Y(_04837_));
 sky130_fd_sc_hd__xnor2_1 _05726_ (.A(_04741_),
    .B(_04826_),
    .Y(_04847_));
 sky130_fd_sc_hd__o21a_1 _05727_ (.A1(_04223_),
    .A2(_04244_),
    .B1(_04847_),
    .X(_04856_));
 sky130_fd_sc_hd__nor3_1 _05728_ (.A(_04223_),
    .B(_04244_),
    .C(_04847_),
    .Y(_04862_));
 sky130_fd_sc_hd__a211oi_2 _05729_ (.A1(_04070_),
    .A2(_04092_),
    .B1(_04856_),
    .C1(_04862_),
    .Y(_04863_));
 sky130_fd_sc_hd__o211a_1 _05730_ (.A1(_04856_),
    .A2(_04862_),
    .B1(_04070_),
    .C1(_04092_),
    .X(_04864_));
 sky130_fd_sc_hd__o21ba_1 _05731_ (.A1(_04179_),
    .A2(_04201_),
    .B1_N(_04168_),
    .X(_04865_));
 sky130_fd_sc_hd__o21ba_1 _05732_ (.A1(_04266_),
    .A2(_04288_),
    .B1_N(_04277_),
    .X(_04866_));
 sky130_fd_sc_hd__and4_1 _05733_ (.A(net471),
    .B(net208),
    .C(net457),
    .D(net199),
    .X(_04867_));
 sky130_fd_sc_hd__a22oi_1 _05734_ (.A1(net208),
    .A2(net457),
    .B1(net199),
    .B2(net471),
    .Y(_04868_));
 sky130_fd_sc_hd__nor2_1 _05735_ (.A(_04867_),
    .B(_04868_),
    .Y(_04869_));
 sky130_fd_sc_hd__nand2_1 _05736_ (.A(net480),
    .B(net196),
    .Y(_04870_));
 sky130_fd_sc_hd__xnor2_1 _05737_ (.A(_04869_),
    .B(_04870_),
    .Y(_04871_));
 sky130_fd_sc_hd__nand2b_1 _05738_ (.A_N(_04866_),
    .B(_04871_),
    .Y(_04872_));
 sky130_fd_sc_hd__xnor2_1 _05739_ (.A(_04866_),
    .B(_04871_),
    .Y(_04873_));
 sky130_fd_sc_hd__nand2b_1 _05740_ (.A_N(_04865_),
    .B(_04873_),
    .Y(_04874_));
 sky130_fd_sc_hd__xnor2_1 _05741_ (.A(_04865_),
    .B(_04873_),
    .Y(_04875_));
 sky130_fd_sc_hd__and4_1 _05742_ (.A(net242),
    .B(net234),
    .C(net546),
    .D(net445),
    .X(_04876_));
 sky130_fd_sc_hd__a22oi_1 _05743_ (.A1(net242),
    .A2(net546),
    .B1(net445),
    .B2(net234),
    .Y(_04877_));
 sky130_fd_sc_hd__nor2_1 _05744_ (.A(_04876_),
    .B(_04877_),
    .Y(_04878_));
 sky130_fd_sc_hd__nand2_1 _05745_ (.A(net217),
    .B(net451),
    .Y(_04879_));
 sky130_fd_sc_hd__xnor2_1 _05746_ (.A(_04878_),
    .B(_04879_),
    .Y(_04880_));
 sky130_fd_sc_hd__nand2_1 _05747_ (.A(net256),
    .B(net465),
    .Y(_04881_));
 sky130_fd_sc_hd__and4_1 _05748_ (.A(net440),
    .B(net347),
    .C(net384),
    .D(net302),
    .X(_04882_));
 sky130_fd_sc_hd__a22oi_2 _05749_ (.A1(net347),
    .A2(net384),
    .B1(net302),
    .B2(net440),
    .Y(_04883_));
 sky130_fd_sc_hd__or3_1 _05750_ (.A(_04881_),
    .B(_04882_),
    .C(_04883_),
    .X(_04884_));
 sky130_fd_sc_hd__o21ai_1 _05751_ (.A1(_04882_),
    .A2(_04883_),
    .B1(_04881_),
    .Y(_04885_));
 sky130_fd_sc_hd__o21bai_1 _05752_ (.A1(_04320_),
    .A2(_04342_),
    .B1_N(_04331_),
    .Y(_04886_));
 sky130_fd_sc_hd__nand3_1 _05753_ (.A(_04884_),
    .B(_04885_),
    .C(_04886_),
    .Y(_04887_));
 sky130_fd_sc_hd__a21o_1 _05754_ (.A1(_04884_),
    .A2(_04885_),
    .B1(_04886_),
    .X(_04888_));
 sky130_fd_sc_hd__nand3_1 _05755_ (.A(_04880_),
    .B(_04887_),
    .C(_04888_),
    .Y(_04889_));
 sky130_fd_sc_hd__a21o_1 _05756_ (.A1(_04887_),
    .A2(_04888_),
    .B1(_04880_),
    .X(_04890_));
 sky130_fd_sc_hd__a21bo_1 _05757_ (.A1(_04310_),
    .A2(_04396_),
    .B1_N(_04385_),
    .X(_04891_));
 sky130_fd_sc_hd__nand3_2 _05758_ (.A(_04889_),
    .B(_04890_),
    .C(_04891_),
    .Y(_04892_));
 sky130_fd_sc_hd__a21o_1 _05759_ (.A1(_04889_),
    .A2(_04890_),
    .B1(_04891_),
    .X(_04893_));
 sky130_fd_sc_hd__and3_1 _05760_ (.A(_04875_),
    .B(_04892_),
    .C(_04893_),
    .X(_04894_));
 sky130_fd_sc_hd__nand3_1 _05761_ (.A(_04875_),
    .B(_04892_),
    .C(_04893_),
    .Y(_04895_));
 sky130_fd_sc_hd__a21oi_1 _05762_ (.A1(_04892_),
    .A2(_04893_),
    .B1(_04875_),
    .Y(_04896_));
 sky130_fd_sc_hd__a211o_1 _05763_ (.A1(_04440_),
    .A2(_04461_),
    .B1(_04894_),
    .C1(_04896_),
    .X(_04897_));
 sky130_fd_sc_hd__o211ai_1 _05764_ (.A1(_04894_),
    .A2(_04896_),
    .B1(_04440_),
    .C1(_04461_),
    .Y(_04898_));
 sky130_fd_sc_hd__or4bb_1 _05765_ (.A(_04863_),
    .B(_04864_),
    .C_N(_04897_),
    .D_N(_04898_),
    .X(_04899_));
 sky130_fd_sc_hd__a2bb2o_1 _05766_ (.A1_N(_04863_),
    .A2_N(_04864_),
    .B1(_04897_),
    .B2(_04898_),
    .X(_04900_));
 sky130_fd_sc_hd__o21bai_1 _05767_ (.A1(_04136_),
    .A2(_04494_),
    .B1_N(_04483_),
    .Y(_04901_));
 sky130_fd_sc_hd__and3_1 _05768_ (.A(_04899_),
    .B(_04900_),
    .C(_04901_),
    .X(_04902_));
 sky130_fd_sc_hd__a21oi_1 _05769_ (.A1(_04899_),
    .A2(_04900_),
    .B1(_04901_),
    .Y(_04903_));
 sky130_fd_sc_hd__nor3_1 _05770_ (.A(_04709_),
    .B(_04902_),
    .C(_04903_),
    .Y(_04904_));
 sky130_fd_sc_hd__o21a_1 _05771_ (.A1(_04902_),
    .A2(_04903_),
    .B1(_04709_),
    .X(_04905_));
 sky130_fd_sc_hd__a21o_1 _05772_ (.A1(_03395_),
    .A2(_04548_),
    .B1(_04537_),
    .X(_04906_));
 sky130_fd_sc_hd__nor3b_1 _05773_ (.A(_04904_),
    .B(_04905_),
    .C_N(_04906_),
    .Y(_04907_));
 sky130_fd_sc_hd__inv_2 _05774_ (.A(_04907_),
    .Y(_04908_));
 sky130_fd_sc_hd__o21ba_1 _05775_ (.A1(_04904_),
    .A2(_04905_),
    .B1_N(_04906_),
    .X(_04909_));
 sky130_fd_sc_hd__nor2_1 _05776_ (.A(_04907_),
    .B(_04909_),
    .Y(_04910_));
 sky130_fd_sc_hd__nand2_1 _05777_ (.A(_04581_),
    .B(_04910_),
    .Y(_04911_));
 sky130_fd_sc_hd__xnor2_2 _05778_ (.A(_04581_),
    .B(_04910_),
    .Y(_04912_));
 sky130_fd_sc_hd__nand3_1 _05779_ (.A(_04602_),
    .B(_04624_),
    .C(_04912_),
    .Y(_04913_));
 sky130_fd_sc_hd__or2_1 _05780_ (.A(_04602_),
    .B(_04912_),
    .X(_04914_));
 sky130_fd_sc_hd__o211ai_2 _05781_ (.A1(_04624_),
    .A2(_04912_),
    .B1(_04913_),
    .C1(_04914_),
    .Y(_04915_));
 sky130_fd_sc_hd__xor2_1 _05782_ (.A(_04698_),
    .B(_04915_),
    .X(net69));
 sky130_fd_sc_hd__o22ai_2 _05783_ (.A1(_04624_),
    .A2(_04912_),
    .B1(_04915_),
    .B2(_04698_),
    .Y(_04916_));
 sky130_fd_sc_hd__o21ai_2 _05784_ (.A1(_04856_),
    .A2(_04863_),
    .B1(_04730_),
    .Y(_04917_));
 sky130_fd_sc_hd__or3_1 _05785_ (.A(_04730_),
    .B(_04856_),
    .C(_04863_),
    .X(_04918_));
 sky130_fd_sc_hd__and2_1 _05786_ (.A(_04917_),
    .B(_04918_),
    .X(_04919_));
 sky130_fd_sc_hd__nand2_1 _05787_ (.A(_04816_),
    .B(_04837_),
    .Y(_04920_));
 sky130_fd_sc_hd__and4_1 _05788_ (.A(net516),
    .B(net600),
    .C(net419),
    .D(net411),
    .X(_04921_));
 sky130_fd_sc_hd__a22oi_1 _05789_ (.A1(net516),
    .A2(net419),
    .B1(net411),
    .B2(net600),
    .Y(_04922_));
 sky130_fd_sc_hd__nor2_1 _05790_ (.A(_04921_),
    .B(_04922_),
    .Y(_04923_));
 sky130_fd_sc_hd__nand2_1 _05791_ (.A(net626),
    .B(net403),
    .Y(_04924_));
 sky130_fd_sc_hd__xnor2_1 _05792_ (.A(_04923_),
    .B(_04924_),
    .Y(_04925_));
 sky130_fd_sc_hd__and4_1 _05793_ (.A(net480),
    .B(net487),
    .C(net191),
    .D(net430),
    .X(_04926_));
 sky130_fd_sc_hd__a22oi_1 _05794_ (.A1(net480),
    .A2(net191),
    .B1(net430),
    .B2(net487),
    .Y(_04927_));
 sky130_fd_sc_hd__nor2_1 _05795_ (.A(_04926_),
    .B(_04927_),
    .Y(_04928_));
 sky130_fd_sc_hd__nand2_1 _05796_ (.A(net495),
    .B(net423),
    .Y(_04929_));
 sky130_fd_sc_hd__xnor2_1 _05797_ (.A(_04928_),
    .B(_04929_),
    .Y(_04930_));
 sky130_fd_sc_hd__o21ba_1 _05798_ (.A1(_04763_),
    .A2(_04784_),
    .B1_N(_04752_),
    .X(_04931_));
 sky130_fd_sc_hd__and2b_1 _05799_ (.A_N(_04931_),
    .B(_04930_),
    .X(_04932_));
 sky130_fd_sc_hd__xnor2_1 _05800_ (.A(_04930_),
    .B(_04931_),
    .Y(_04933_));
 sky130_fd_sc_hd__and2_1 _05801_ (.A(_04925_),
    .B(_04933_),
    .X(_04934_));
 sky130_fd_sc_hd__xnor2_1 _05802_ (.A(_04925_),
    .B(_04933_),
    .Y(_04935_));
 sky130_fd_sc_hd__a21o_1 _05803_ (.A1(_04872_),
    .A2(_04874_),
    .B1(_04935_),
    .X(_04936_));
 sky130_fd_sc_hd__nand3_1 _05804_ (.A(_04872_),
    .B(_04874_),
    .C(_04935_),
    .Y(_04937_));
 sky130_fd_sc_hd__nand3_1 _05805_ (.A(_04920_),
    .B(_04936_),
    .C(_04937_),
    .Y(_04938_));
 sky130_fd_sc_hd__a21o_1 _05806_ (.A1(_04936_),
    .A2(_04937_),
    .B1(_04920_),
    .X(_04939_));
 sky130_fd_sc_hd__o21ba_1 _05807_ (.A1(_04868_),
    .A2(_04870_),
    .B1_N(_04867_),
    .X(_04940_));
 sky130_fd_sc_hd__o21ba_1 _05808_ (.A1(_04877_),
    .A2(_04879_),
    .B1_N(_04876_),
    .X(_04941_));
 sky130_fd_sc_hd__and4_1 _05809_ (.A(net214),
    .B(net457),
    .C(net199),
    .D(net452),
    .X(_04942_));
 sky130_fd_sc_hd__a22oi_1 _05810_ (.A1(net457),
    .A2(net199),
    .B1(net452),
    .B2(net214),
    .Y(_04943_));
 sky130_fd_sc_hd__nor2_1 _05811_ (.A(_04942_),
    .B(_04943_),
    .Y(_04944_));
 sky130_fd_sc_hd__nand2_1 _05812_ (.A(net472),
    .B(net196),
    .Y(_04945_));
 sky130_fd_sc_hd__xnor2_1 _05813_ (.A(_04944_),
    .B(_04945_),
    .Y(_04946_));
 sky130_fd_sc_hd__nand2b_1 _05814_ (.A_N(_04941_),
    .B(_04946_),
    .Y(_04947_));
 sky130_fd_sc_hd__xnor2_1 _05815_ (.A(_04941_),
    .B(_04946_),
    .Y(_04948_));
 sky130_fd_sc_hd__nand2b_1 _05816_ (.A_N(_04940_),
    .B(_04948_),
    .Y(_04949_));
 sky130_fd_sc_hd__xnor2_1 _05817_ (.A(_04940_),
    .B(_04948_),
    .Y(_04950_));
 sky130_fd_sc_hd__and4_1 _05818_ (.A(net242),
    .B(net234),
    .C(net546),
    .D(net465),
    .X(_04951_));
 sky130_fd_sc_hd__a22oi_1 _05819_ (.A1(net234),
    .A2(net546),
    .B1(net465),
    .B2(net242),
    .Y(_04952_));
 sky130_fd_sc_hd__nor2_1 _05820_ (.A(_04951_),
    .B(_04952_),
    .Y(_04953_));
 sky130_fd_sc_hd__nand2_1 _05821_ (.A(net217),
    .B(net445),
    .Y(_04954_));
 sky130_fd_sc_hd__xnor2_1 _05822_ (.A(_04953_),
    .B(_04954_),
    .Y(_04955_));
 sky130_fd_sc_hd__nand2_1 _05823_ (.A(net256),
    .B(net384),
    .Y(_04956_));
 sky130_fd_sc_hd__and4_1 _05824_ (.A(net440),
    .B(net347),
    .C(net302),
    .D(net226),
    .X(_04957_));
 sky130_fd_sc_hd__a22oi_2 _05825_ (.A1(net347),
    .A2(net302),
    .B1(net226),
    .B2(net440),
    .Y(_04958_));
 sky130_fd_sc_hd__or3_1 _05826_ (.A(_04956_),
    .B(_04957_),
    .C(_04958_),
    .X(_04959_));
 sky130_fd_sc_hd__o21ai_1 _05827_ (.A1(_04957_),
    .A2(_04958_),
    .B1(_04956_),
    .Y(_04960_));
 sky130_fd_sc_hd__o21bai_1 _05828_ (.A1(_04881_),
    .A2(_04883_),
    .B1_N(_04882_),
    .Y(_04961_));
 sky130_fd_sc_hd__nand3_1 _05829_ (.A(_04959_),
    .B(_04960_),
    .C(_04961_),
    .Y(_04962_));
 sky130_fd_sc_hd__a21o_1 _05830_ (.A1(_04959_),
    .A2(_04960_),
    .B1(_04961_),
    .X(_04963_));
 sky130_fd_sc_hd__nand3_1 _05831_ (.A(_04955_),
    .B(_04962_),
    .C(_04963_),
    .Y(_04964_));
 sky130_fd_sc_hd__a21o_1 _05832_ (.A1(_04962_),
    .A2(_04963_),
    .B1(_04955_),
    .X(_04965_));
 sky130_fd_sc_hd__a21bo_1 _05833_ (.A1(_04880_),
    .A2(_04888_),
    .B1_N(_04887_),
    .X(_04966_));
 sky130_fd_sc_hd__nand3_2 _05834_ (.A(_04964_),
    .B(_04965_),
    .C(_04966_),
    .Y(_04967_));
 sky130_fd_sc_hd__a21o_1 _05835_ (.A1(_04964_),
    .A2(_04965_),
    .B1(_04966_),
    .X(_04968_));
 sky130_fd_sc_hd__and3_1 _05836_ (.A(_04950_),
    .B(_04967_),
    .C(_04968_),
    .X(_04969_));
 sky130_fd_sc_hd__nand3_1 _05837_ (.A(_04950_),
    .B(_04967_),
    .C(_04968_),
    .Y(_04970_));
 sky130_fd_sc_hd__a21oi_1 _05838_ (.A1(_04967_),
    .A2(_04968_),
    .B1(_04950_),
    .Y(_04971_));
 sky130_fd_sc_hd__a211o_1 _05839_ (.A1(_04892_),
    .A2(_04895_),
    .B1(_04969_),
    .C1(_04971_),
    .X(_04972_));
 sky130_fd_sc_hd__o211ai_2 _05840_ (.A1(_04969_),
    .A2(_04971_),
    .B1(_04892_),
    .C1(_04895_),
    .Y(_04973_));
 sky130_fd_sc_hd__and4_1 _05841_ (.A(_04938_),
    .B(_04939_),
    .C(_04972_),
    .D(_04973_),
    .X(_04974_));
 sky130_fd_sc_hd__nand4_1 _05842_ (.A(_04938_),
    .B(_04939_),
    .C(_04972_),
    .D(_04973_),
    .Y(_04975_));
 sky130_fd_sc_hd__a22oi_1 _05843_ (.A1(_04938_),
    .A2(_04939_),
    .B1(_04972_),
    .B2(_04973_),
    .Y(_04976_));
 sky130_fd_sc_hd__a211o_1 _05844_ (.A1(_04897_),
    .A2(_04899_),
    .B1(_04974_),
    .C1(_04976_),
    .X(_04977_));
 sky130_fd_sc_hd__o211ai_1 _05845_ (.A1(_04974_),
    .A2(_04976_),
    .B1(_04897_),
    .C1(_04899_),
    .Y(_04978_));
 sky130_fd_sc_hd__nand3_1 _05846_ (.A(_04919_),
    .B(_04977_),
    .C(_04978_),
    .Y(_04979_));
 sky130_fd_sc_hd__a21o_1 _05847_ (.A1(_04977_),
    .A2(_04978_),
    .B1(_04919_),
    .X(_04980_));
 sky130_fd_sc_hd__nand2_1 _05848_ (.A(_04979_),
    .B(_04980_),
    .Y(_04981_));
 sky130_fd_sc_hd__nor2_1 _05849_ (.A(_04902_),
    .B(_04904_),
    .Y(_04982_));
 sky130_fd_sc_hd__nor2_2 _05850_ (.A(_04981_),
    .B(_04982_),
    .Y(_04983_));
 sky130_fd_sc_hd__xnor2_1 _05851_ (.A(_04981_),
    .B(_04982_),
    .Y(_04984_));
 sky130_fd_sc_hd__or2_1 _05852_ (.A(_04908_),
    .B(_04984_),
    .X(_04985_));
 sky130_fd_sc_hd__nand2_1 _05853_ (.A(_04908_),
    .B(_04984_),
    .Y(_04986_));
 sky130_fd_sc_hd__nand2_1 _05854_ (.A(_04985_),
    .B(_04986_),
    .Y(_04987_));
 sky130_fd_sc_hd__nor2_1 _05855_ (.A(_04911_),
    .B(_04987_),
    .Y(_04988_));
 sky130_fd_sc_hd__nand2_1 _05856_ (.A(_04911_),
    .B(_04914_),
    .Y(_04989_));
 sky130_fd_sc_hd__xnor2_1 _05857_ (.A(_04987_),
    .B(_04989_),
    .Y(_04990_));
 sky130_fd_sc_hd__xor2_1 _05858_ (.A(_04916_),
    .B(_04990_),
    .X(net70));
 sky130_fd_sc_hd__a2bb2o_1 _05859_ (.A1_N(_04914_),
    .A2_N(_04987_),
    .B1(_04990_),
    .B2(_04916_),
    .X(_04991_));
 sky130_fd_sc_hd__o21ba_1 _05860_ (.A1(_04922_),
    .A2(_04924_),
    .B1_N(_04921_),
    .X(_04992_));
 sky130_fd_sc_hd__nand2_1 _05861_ (.A(net626),
    .B(net396),
    .Y(_04993_));
 sky130_fd_sc_hd__nor2_1 _05862_ (.A(_04992_),
    .B(_04993_),
    .Y(_04994_));
 sky130_fd_sc_hd__xnor2_1 _05863_ (.A(_04992_),
    .B(_04993_),
    .Y(_04995_));
 sky130_fd_sc_hd__a21oi_1 _05864_ (.A1(_04936_),
    .A2(_04938_),
    .B1(_04995_),
    .Y(_04996_));
 sky130_fd_sc_hd__and3_1 _05865_ (.A(_04936_),
    .B(_04938_),
    .C(_04995_),
    .X(_04997_));
 sky130_fd_sc_hd__nor2_1 _05866_ (.A(_04996_),
    .B(_04997_),
    .Y(_04998_));
 sky130_fd_sc_hd__and4_1 _05867_ (.A(net495),
    .B(net516),
    .C(net419),
    .D(net411),
    .X(_04999_));
 sky130_fd_sc_hd__a22oi_1 _05868_ (.A1(net495),
    .A2(net419),
    .B1(net411),
    .B2(net516),
    .Y(_05000_));
 sky130_fd_sc_hd__nor2_1 _05869_ (.A(_04999_),
    .B(_05000_),
    .Y(_05001_));
 sky130_fd_sc_hd__a21oi_1 _05870_ (.A1(net600),
    .A2(net403),
    .B1(_05001_),
    .Y(_05002_));
 sky130_fd_sc_hd__and3_1 _05871_ (.A(net600),
    .B(net403),
    .C(_05001_),
    .X(_05003_));
 sky130_fd_sc_hd__nor2_1 _05872_ (.A(_05002_),
    .B(_05003_),
    .Y(_05004_));
 sky130_fd_sc_hd__and4_1 _05873_ (.A(net480),
    .B(net472),
    .C(net188),
    .D(net433),
    .X(_05005_));
 sky130_fd_sc_hd__a22o_1 _05874_ (.A1(net472),
    .A2(net188),
    .B1(net433),
    .B2(net480),
    .X(_05006_));
 sky130_fd_sc_hd__and2b_1 _05875_ (.A_N(_05005_),
    .B(_05006_),
    .X(_05007_));
 sky130_fd_sc_hd__nand2_1 _05876_ (.A(net487),
    .B(net423),
    .Y(_05008_));
 sky130_fd_sc_hd__xnor2_1 _05877_ (.A(_05007_),
    .B(_05008_),
    .Y(_05009_));
 sky130_fd_sc_hd__o21ba_1 _05878_ (.A1(_04927_),
    .A2(_04929_),
    .B1_N(_04926_),
    .X(_05010_));
 sky130_fd_sc_hd__and2b_1 _05879_ (.A_N(_05010_),
    .B(_05009_),
    .X(_05011_));
 sky130_fd_sc_hd__xnor2_1 _05880_ (.A(_05009_),
    .B(_05010_),
    .Y(_05012_));
 sky130_fd_sc_hd__and2_1 _05881_ (.A(_05004_),
    .B(_05012_),
    .X(_05013_));
 sky130_fd_sc_hd__xnor2_1 _05882_ (.A(_05004_),
    .B(_05012_),
    .Y(_05014_));
 sky130_fd_sc_hd__a21o_1 _05883_ (.A1(_04947_),
    .A2(_04949_),
    .B1(_05014_),
    .X(_05015_));
 sky130_fd_sc_hd__nand3_2 _05884_ (.A(_04947_),
    .B(_04949_),
    .C(_05014_),
    .Y(_05016_));
 sky130_fd_sc_hd__o211ai_4 _05885_ (.A1(_04932_),
    .A2(_04934_),
    .B1(_05015_),
    .C1(_05016_),
    .Y(_05017_));
 sky130_fd_sc_hd__a211o_1 _05886_ (.A1(_05015_),
    .A2(_05016_),
    .B1(_04932_),
    .C1(_04934_),
    .X(_05018_));
 sky130_fd_sc_hd__a31o_1 _05887_ (.A1(net472),
    .A2(net196),
    .A3(_04944_),
    .B1(_04942_),
    .X(_05019_));
 sky130_fd_sc_hd__o21bai_1 _05888_ (.A1(_04952_),
    .A2(_04954_),
    .B1_N(_04951_),
    .Y(_05020_));
 sky130_fd_sc_hd__nand4_1 _05889_ (.A(net214),
    .B(net205),
    .C(net452),
    .D(net446),
    .Y(_05021_));
 sky130_fd_sc_hd__a22o_1 _05890_ (.A1(net205),
    .A2(net452),
    .B1(net446),
    .B2(net214),
    .X(_05022_));
 sky130_fd_sc_hd__a22o_1 _05891_ (.A1(net457),
    .A2(net196),
    .B1(_05021_),
    .B2(_05022_),
    .X(_05023_));
 sky130_fd_sc_hd__nand4_1 _05892_ (.A(net457),
    .B(net196),
    .C(_05021_),
    .D(_05022_),
    .Y(_05024_));
 sky130_fd_sc_hd__and3_1 _05893_ (.A(_05020_),
    .B(_05023_),
    .C(_05024_),
    .X(_05025_));
 sky130_fd_sc_hd__a21o_1 _05894_ (.A1(_05023_),
    .A2(_05024_),
    .B1(_05020_),
    .X(_05026_));
 sky130_fd_sc_hd__and2b_1 _05895_ (.A_N(_05025_),
    .B(_05026_),
    .X(_05027_));
 sky130_fd_sc_hd__xor2_1 _05896_ (.A(_05019_),
    .B(_05027_),
    .X(_05028_));
 sky130_fd_sc_hd__and4_1 _05897_ (.A(net242),
    .B(net234),
    .C(net465),
    .D(net384),
    .X(_05029_));
 sky130_fd_sc_hd__a22oi_1 _05898_ (.A1(net234),
    .A2(net465),
    .B1(net384),
    .B2(net242),
    .Y(_05030_));
 sky130_fd_sc_hd__nor2_1 _05899_ (.A(_05029_),
    .B(_05030_),
    .Y(_05031_));
 sky130_fd_sc_hd__nand2_1 _05900_ (.A(net217),
    .B(net546),
    .Y(_05032_));
 sky130_fd_sc_hd__xnor2_1 _05901_ (.A(_05031_),
    .B(_05032_),
    .Y(_05033_));
 sky130_fd_sc_hd__nand2_1 _05902_ (.A(net256),
    .B(net302),
    .Y(_05034_));
 sky130_fd_sc_hd__and4_1 _05903_ (.A(net440),
    .B(net347),
    .C(net226),
    .D(net181),
    .X(_05035_));
 sky130_fd_sc_hd__a22oi_2 _05904_ (.A1(net347),
    .A2(net226),
    .B1(net181),
    .B2(net440),
    .Y(_05036_));
 sky130_fd_sc_hd__or3_1 _05905_ (.A(_05034_),
    .B(_05035_),
    .C(_05036_),
    .X(_05037_));
 sky130_fd_sc_hd__o21ai_1 _05906_ (.A1(_05035_),
    .A2(_05036_),
    .B1(_05034_),
    .Y(_05038_));
 sky130_fd_sc_hd__o21bai_1 _05907_ (.A1(_04956_),
    .A2(_04958_),
    .B1_N(_04957_),
    .Y(_05039_));
 sky130_fd_sc_hd__nand3_1 _05908_ (.A(_05037_),
    .B(_05038_),
    .C(_05039_),
    .Y(_05040_));
 sky130_fd_sc_hd__a21o_1 _05909_ (.A1(_05037_),
    .A2(_05038_),
    .B1(_05039_),
    .X(_05041_));
 sky130_fd_sc_hd__nand3_1 _05910_ (.A(_05033_),
    .B(_05040_),
    .C(_05041_),
    .Y(_05042_));
 sky130_fd_sc_hd__a21o_1 _05911_ (.A1(_05040_),
    .A2(_05041_),
    .B1(_05033_),
    .X(_05043_));
 sky130_fd_sc_hd__a21bo_1 _05912_ (.A1(_04955_),
    .A2(_04963_),
    .B1_N(_04962_),
    .X(_05044_));
 sky130_fd_sc_hd__nand3_4 _05913_ (.A(_05042_),
    .B(_05043_),
    .C(_05044_),
    .Y(_05045_));
 sky130_fd_sc_hd__a21o_1 _05914_ (.A1(_05042_),
    .A2(_05043_),
    .B1(_05044_),
    .X(_05046_));
 sky130_fd_sc_hd__and3_1 _05915_ (.A(_05028_),
    .B(_05045_),
    .C(_05046_),
    .X(_05047_));
 sky130_fd_sc_hd__nand3_2 _05916_ (.A(_05028_),
    .B(_05045_),
    .C(_05046_),
    .Y(_05048_));
 sky130_fd_sc_hd__a21oi_1 _05917_ (.A1(_05045_),
    .A2(_05046_),
    .B1(_05028_),
    .Y(_05049_));
 sky130_fd_sc_hd__a211o_1 _05918_ (.A1(_04967_),
    .A2(_04970_),
    .B1(_05047_),
    .C1(_05049_),
    .X(_05050_));
 sky130_fd_sc_hd__o211ai_2 _05919_ (.A1(_05047_),
    .A2(_05049_),
    .B1(_04967_),
    .C1(_04970_),
    .Y(_05051_));
 sky130_fd_sc_hd__and4_1 _05920_ (.A(_05017_),
    .B(_05018_),
    .C(_05050_),
    .D(_05051_),
    .X(_05052_));
 sky130_fd_sc_hd__nand4_1 _05921_ (.A(_05017_),
    .B(_05018_),
    .C(_05050_),
    .D(_05051_),
    .Y(_05053_));
 sky130_fd_sc_hd__a22oi_2 _05922_ (.A1(_05017_),
    .A2(_05018_),
    .B1(_05050_),
    .B2(_05051_),
    .Y(_05054_));
 sky130_fd_sc_hd__a211o_1 _05923_ (.A1(_04972_),
    .A2(_04975_),
    .B1(_05052_),
    .C1(_05054_),
    .X(_05055_));
 sky130_fd_sc_hd__inv_2 _05924_ (.A(_05055_),
    .Y(_05056_));
 sky130_fd_sc_hd__o211ai_1 _05925_ (.A1(_05052_),
    .A2(_05054_),
    .B1(_04972_),
    .C1(_04975_),
    .Y(_05057_));
 sky130_fd_sc_hd__and3_1 _05926_ (.A(_04998_),
    .B(_05055_),
    .C(_05057_),
    .X(_05058_));
 sky130_fd_sc_hd__a21oi_1 _05927_ (.A1(_05055_),
    .A2(_05057_),
    .B1(_04998_),
    .Y(_05059_));
 sky130_fd_sc_hd__or2_1 _05928_ (.A(_05058_),
    .B(_05059_),
    .X(_05060_));
 sky130_fd_sc_hd__nand2_1 _05929_ (.A(_04977_),
    .B(_04979_),
    .Y(_05061_));
 sky130_fd_sc_hd__a211oi_1 _05930_ (.A1(_04977_),
    .A2(_04979_),
    .B1(_05058_),
    .C1(_05059_),
    .Y(_05062_));
 sky130_fd_sc_hd__xnor2_1 _05931_ (.A(_05060_),
    .B(_05061_),
    .Y(_05063_));
 sky130_fd_sc_hd__a211oi_1 _05932_ (.A1(_04977_),
    .A2(_05060_),
    .B1(_05062_),
    .C1(_04917_),
    .Y(_05064_));
 sky130_fd_sc_hd__xnor2_2 _05933_ (.A(_04917_),
    .B(_05063_),
    .Y(_05065_));
 sky130_fd_sc_hd__and2_1 _05934_ (.A(_04983_),
    .B(_05065_),
    .X(_05066_));
 sky130_fd_sc_hd__xor2_4 _05935_ (.A(_04983_),
    .B(_05065_),
    .X(_05067_));
 sky130_fd_sc_hd__o21a_1 _05936_ (.A1(_04911_),
    .A2(_04987_),
    .B1(_04985_),
    .X(_05068_));
 sky130_fd_sc_hd__xnor2_2 _05937_ (.A(_05067_),
    .B(_05068_),
    .Y(_05069_));
 sky130_fd_sc_hd__xor2_1 _05938_ (.A(_04991_),
    .B(_05069_),
    .X(net71));
 sky130_fd_sc_hd__a22oi_4 _05939_ (.A1(_04988_),
    .A2(_05067_),
    .B1(_05069_),
    .B2(_04991_),
    .Y(_05070_));
 sky130_fd_sc_hd__nand2b_1 _05940_ (.A_N(_04985_),
    .B(_05067_),
    .Y(_05071_));
 sky130_fd_sc_hd__and4_1 _05941_ (.A(net600),
    .B(net626),
    .C(net396),
    .D(net380),
    .X(_05072_));
 sky130_fd_sc_hd__nand4_1 _05942_ (.A(net601),
    .B(net626),
    .C(net396),
    .D(net380),
    .Y(_05073_));
 sky130_fd_sc_hd__a22o_1 _05943_ (.A1(net601),
    .A2(net396),
    .B1(net380),
    .B2(net626),
    .X(_05074_));
 sky130_fd_sc_hd__o211a_1 _05944_ (.A1(_04999_),
    .A2(_05003_),
    .B1(_05073_),
    .C1(_05074_),
    .X(_05075_));
 sky130_fd_sc_hd__a211oi_1 _05945_ (.A1(_05073_),
    .A2(_05074_),
    .B1(_04999_),
    .C1(_05003_),
    .Y(_05076_));
 sky130_fd_sc_hd__nor2_1 _05946_ (.A(_05075_),
    .B(_05076_),
    .Y(_05077_));
 sky130_fd_sc_hd__nand2_1 _05947_ (.A(_04994_),
    .B(_05077_),
    .Y(_05078_));
 sky130_fd_sc_hd__or2_1 _05948_ (.A(_04994_),
    .B(_05077_),
    .X(_05079_));
 sky130_fd_sc_hd__nand2_1 _05949_ (.A(_05078_),
    .B(_05079_),
    .Y(_05080_));
 sky130_fd_sc_hd__a21oi_1 _05950_ (.A1(_05015_),
    .A2(_05017_),
    .B1(_05080_),
    .Y(_05081_));
 sky130_fd_sc_hd__and3_1 _05951_ (.A(_05015_),
    .B(_05017_),
    .C(_05080_),
    .X(_05082_));
 sky130_fd_sc_hd__nor2_1 _05952_ (.A(_05081_),
    .B(_05082_),
    .Y(_05083_));
 sky130_fd_sc_hd__a21o_1 _05953_ (.A1(_05019_),
    .A2(_05026_),
    .B1(_05025_),
    .X(_05084_));
 sky130_fd_sc_hd__and4_1 _05954_ (.A(net487),
    .B(net495),
    .C(net419),
    .D(net411),
    .X(_05085_));
 sky130_fd_sc_hd__a22o_1 _05955_ (.A1(net487),
    .A2(net419),
    .B1(net411),
    .B2(net495),
    .X(_05086_));
 sky130_fd_sc_hd__and2b_1 _05956_ (.A_N(_05085_),
    .B(_05086_),
    .X(_05087_));
 sky130_fd_sc_hd__nand2_1 _05957_ (.A(net516),
    .B(net403),
    .Y(_05088_));
 sky130_fd_sc_hd__xnor2_1 _05958_ (.A(_05087_),
    .B(_05088_),
    .Y(_05089_));
 sky130_fd_sc_hd__nand4_1 _05959_ (.A(net472),
    .B(net457),
    .C(net188),
    .D(net431),
    .Y(_05090_));
 sky130_fd_sc_hd__a22o_1 _05960_ (.A1(net457),
    .A2(net188),
    .B1(net431),
    .B2(net472),
    .X(_05091_));
 sky130_fd_sc_hd__and2_1 _05961_ (.A(net480),
    .B(net423),
    .X(_05092_));
 sky130_fd_sc_hd__a21o_1 _05962_ (.A1(_05090_),
    .A2(_05091_),
    .B1(_05092_),
    .X(_05093_));
 sky130_fd_sc_hd__nand3_1 _05963_ (.A(_05090_),
    .B(_05091_),
    .C(_05092_),
    .Y(_05094_));
 sky130_fd_sc_hd__a31o_1 _05964_ (.A1(net487),
    .A2(net423),
    .A3(_05006_),
    .B1(_05005_),
    .X(_05095_));
 sky130_fd_sc_hd__nand3_1 _05965_ (.A(_05093_),
    .B(_05094_),
    .C(_05095_),
    .Y(_05096_));
 sky130_fd_sc_hd__a21o_1 _05966_ (.A1(_05093_),
    .A2(_05094_),
    .B1(_05095_),
    .X(_05097_));
 sky130_fd_sc_hd__nand3_1 _05967_ (.A(_05089_),
    .B(_05096_),
    .C(_05097_),
    .Y(_05098_));
 sky130_fd_sc_hd__a21o_1 _05968_ (.A1(_05096_),
    .A2(_05097_),
    .B1(_05089_),
    .X(_05099_));
 sky130_fd_sc_hd__nand3_2 _05969_ (.A(_05084_),
    .B(_05098_),
    .C(_05099_),
    .Y(_05100_));
 sky130_fd_sc_hd__a21o_1 _05970_ (.A1(_05098_),
    .A2(_05099_),
    .B1(_05084_),
    .X(_05101_));
 sky130_fd_sc_hd__o211ai_2 _05971_ (.A1(_05011_),
    .A2(_05013_),
    .B1(_05100_),
    .C1(_05101_),
    .Y(_05102_));
 sky130_fd_sc_hd__a211o_1 _05972_ (.A1(_05100_),
    .A2(_05101_),
    .B1(_05011_),
    .C1(_05013_),
    .X(_05103_));
 sky130_fd_sc_hd__nand2_1 _05973_ (.A(_05102_),
    .B(_05103_),
    .Y(_05104_));
 sky130_fd_sc_hd__nand2_1 _05974_ (.A(_05021_),
    .B(_05024_),
    .Y(_05105_));
 sky130_fd_sc_hd__o21bai_1 _05975_ (.A1(_05030_),
    .A2(_05032_),
    .B1_N(_05029_),
    .Y(_05106_));
 sky130_fd_sc_hd__nand4_1 _05976_ (.A(net214),
    .B(net205),
    .C(net547),
    .D(net446),
    .Y(_05107_));
 sky130_fd_sc_hd__a22o_1 _05977_ (.A1(net214),
    .A2(net547),
    .B1(net446),
    .B2(net205),
    .X(_05108_));
 sky130_fd_sc_hd__a22o_1 _05978_ (.A1(net452),
    .A2(net195),
    .B1(_05107_),
    .B2(_05108_),
    .X(_05109_));
 sky130_fd_sc_hd__nand4_1 _05979_ (.A(net452),
    .B(net195),
    .C(_05107_),
    .D(_05108_),
    .Y(_05110_));
 sky130_fd_sc_hd__and3_1 _05980_ (.A(_05106_),
    .B(_05109_),
    .C(_05110_),
    .X(_05111_));
 sky130_fd_sc_hd__a21o_1 _05981_ (.A1(_05109_),
    .A2(_05110_),
    .B1(_05106_),
    .X(_05112_));
 sky130_fd_sc_hd__and2b_1 _05982_ (.A_N(_05111_),
    .B(_05112_),
    .X(_05113_));
 sky130_fd_sc_hd__xor2_1 _05983_ (.A(_05105_),
    .B(_05113_),
    .X(_05114_));
 sky130_fd_sc_hd__and4_1 _05984_ (.A(net240),
    .B(net232),
    .C(net384),
    .D(net302),
    .X(_05115_));
 sky130_fd_sc_hd__a22oi_1 _05985_ (.A1(net232),
    .A2(net384),
    .B1(net302),
    .B2(net240),
    .Y(_05116_));
 sky130_fd_sc_hd__nor2_1 _05986_ (.A(_05115_),
    .B(_05116_),
    .Y(_05117_));
 sky130_fd_sc_hd__nand2_1 _05987_ (.A(net217),
    .B(net465),
    .Y(_05118_));
 sky130_fd_sc_hd__xnor2_1 _05988_ (.A(_05117_),
    .B(_05118_),
    .Y(_05119_));
 sky130_fd_sc_hd__nand2_1 _05989_ (.A(net256),
    .B(net226),
    .Y(_05120_));
 sky130_fd_sc_hd__and4_1 _05990_ (.A(net439),
    .B(net346),
    .C(net181),
    .D(net174),
    .X(_05121_));
 sky130_fd_sc_hd__a22oi_2 _05991_ (.A1(net346),
    .A2(net181),
    .B1(net174),
    .B2(net439),
    .Y(_05122_));
 sky130_fd_sc_hd__or3_1 _05992_ (.A(_05120_),
    .B(_05121_),
    .C(_05122_),
    .X(_05123_));
 sky130_fd_sc_hd__o21ai_1 _05993_ (.A1(_05121_),
    .A2(_05122_),
    .B1(_05120_),
    .Y(_05124_));
 sky130_fd_sc_hd__o21bai_1 _05994_ (.A1(_05034_),
    .A2(_05036_),
    .B1_N(_05035_),
    .Y(_05125_));
 sky130_fd_sc_hd__nand3_1 _05995_ (.A(_05123_),
    .B(_05124_),
    .C(_05125_),
    .Y(_05126_));
 sky130_fd_sc_hd__a21o_1 _05996_ (.A1(_05123_),
    .A2(_05124_),
    .B1(_05125_),
    .X(_05127_));
 sky130_fd_sc_hd__nand3_1 _05997_ (.A(_05119_),
    .B(_05126_),
    .C(_05127_),
    .Y(_05128_));
 sky130_fd_sc_hd__a21o_1 _05998_ (.A1(_05126_),
    .A2(_05127_),
    .B1(_05119_),
    .X(_05129_));
 sky130_fd_sc_hd__a21bo_1 _05999_ (.A1(_05033_),
    .A2(_05041_),
    .B1_N(_05040_),
    .X(_05130_));
 sky130_fd_sc_hd__nand3_2 _06000_ (.A(_05128_),
    .B(_05129_),
    .C(_05130_),
    .Y(_05131_));
 sky130_fd_sc_hd__a21o_1 _06001_ (.A1(_05128_),
    .A2(_05129_),
    .B1(_05130_),
    .X(_05132_));
 sky130_fd_sc_hd__and3_1 _06002_ (.A(_05114_),
    .B(_05131_),
    .C(_05132_),
    .X(_05133_));
 sky130_fd_sc_hd__nand3_1 _06003_ (.A(_05114_),
    .B(_05131_),
    .C(_05132_),
    .Y(_05134_));
 sky130_fd_sc_hd__a21oi_2 _06004_ (.A1(_05131_),
    .A2(_05132_),
    .B1(_05114_),
    .Y(_05135_));
 sky130_fd_sc_hd__a211oi_4 _06005_ (.A1(_05045_),
    .A2(_05048_),
    .B1(_05133_),
    .C1(_05135_),
    .Y(_05136_));
 sky130_fd_sc_hd__o211a_1 _06006_ (.A1(_05133_),
    .A2(_05135_),
    .B1(_05045_),
    .C1(_05048_),
    .X(_05137_));
 sky130_fd_sc_hd__nor3_2 _06007_ (.A(_05104_),
    .B(_05136_),
    .C(_05137_),
    .Y(_05138_));
 sky130_fd_sc_hd__o21a_1 _06008_ (.A1(_05136_),
    .A2(_05137_),
    .B1(_05104_),
    .X(_05139_));
 sky130_fd_sc_hd__a211o_1 _06009_ (.A1(_05050_),
    .A2(_05053_),
    .B1(_05138_),
    .C1(_05139_),
    .X(_05140_));
 sky130_fd_sc_hd__o211ai_2 _06010_ (.A1(_05138_),
    .A2(_05139_),
    .B1(_05050_),
    .C1(_05053_),
    .Y(_05141_));
 sky130_fd_sc_hd__nand3_2 _06011_ (.A(_05083_),
    .B(_05140_),
    .C(_05141_),
    .Y(_05142_));
 sky130_fd_sc_hd__a21o_1 _06012_ (.A1(_05140_),
    .A2(_05141_),
    .B1(_05083_),
    .X(_05143_));
 sky130_fd_sc_hd__o211ai_2 _06013_ (.A1(_05056_),
    .A2(_05058_),
    .B1(_05142_),
    .C1(_05143_),
    .Y(_05144_));
 sky130_fd_sc_hd__a211o_1 _06014_ (.A1(_05142_),
    .A2(_05143_),
    .B1(_05056_),
    .C1(_05058_),
    .X(_05145_));
 sky130_fd_sc_hd__nand3_1 _06015_ (.A(_04996_),
    .B(_05144_),
    .C(_05145_),
    .Y(_05146_));
 sky130_fd_sc_hd__a21o_1 _06016_ (.A1(_05144_),
    .A2(_05145_),
    .B1(_04996_),
    .X(_05147_));
 sky130_fd_sc_hd__o211a_1 _06017_ (.A1(_05062_),
    .A2(_05064_),
    .B1(_05146_),
    .C1(_05147_),
    .X(_05148_));
 sky130_fd_sc_hd__a211oi_1 _06018_ (.A1(_05146_),
    .A2(_05147_),
    .B1(_05062_),
    .C1(_05064_),
    .Y(_05149_));
 sky130_fd_sc_hd__nor2_1 _06019_ (.A(_05148_),
    .B(_05149_),
    .Y(_05150_));
 sky130_fd_sc_hd__nor2_1 _06020_ (.A(_05066_),
    .B(_05150_),
    .Y(_05151_));
 sky130_fd_sc_hd__nand2_1 _06021_ (.A(_05071_),
    .B(_05151_),
    .Y(_05152_));
 sky130_fd_sc_hd__nand2_1 _06022_ (.A(_05066_),
    .B(_05150_),
    .Y(_05153_));
 sky130_fd_sc_hd__o311a_1 _06023_ (.A1(_05071_),
    .A2(_05148_),
    .A3(_05149_),
    .B1(_05152_),
    .C1(_05153_),
    .X(_05154_));
 sky130_fd_sc_hd__nand2b_1 _06024_ (.A_N(_05070_),
    .B(_05154_),
    .Y(_05155_));
 sky130_fd_sc_hd__xnor2_1 _06025_ (.A(_05070_),
    .B(_05154_),
    .Y(net72));
 sky130_fd_sc_hd__o31a_1 _06026_ (.A1(_05071_),
    .A2(_05148_),
    .A3(_05149_),
    .B1(_05155_),
    .X(_05156_));
 sky130_fd_sc_hd__a31o_1 _06027_ (.A1(net516),
    .A2(net403),
    .A3(_05086_),
    .B1(_05085_),
    .X(_05157_));
 sky130_fd_sc_hd__and4_1 _06028_ (.A(net516),
    .B(net604),
    .C(net396),
    .D(net380),
    .X(_05158_));
 sky130_fd_sc_hd__a22oi_1 _06029_ (.A1(net520),
    .A2(net396),
    .B1(net380),
    .B2(net601),
    .Y(_05159_));
 sky130_fd_sc_hd__and4bb_1 _06030_ (.A_N(_05158_),
    .B_N(_05159_),
    .C(net629),
    .D(net372),
    .X(_05160_));
 sky130_fd_sc_hd__o2bb2a_1 _06031_ (.A1_N(net629),
    .A2_N(net372),
    .B1(_05158_),
    .B2(_05159_),
    .X(_05161_));
 sky130_fd_sc_hd__nor2_1 _06032_ (.A(_05160_),
    .B(_05161_),
    .Y(_05162_));
 sky130_fd_sc_hd__or2_1 _06033_ (.A(_05157_),
    .B(_05162_),
    .X(_05163_));
 sky130_fd_sc_hd__and2_1 _06034_ (.A(_05157_),
    .B(_05162_),
    .X(_05164_));
 sky130_fd_sc_hd__nand2_1 _06035_ (.A(_05157_),
    .B(_05162_),
    .Y(_05165_));
 sky130_fd_sc_hd__nand2_1 _06036_ (.A(_05163_),
    .B(_05165_),
    .Y(_05166_));
 sky130_fd_sc_hd__nor2_1 _06037_ (.A(_05072_),
    .B(_05075_),
    .Y(_05167_));
 sky130_fd_sc_hd__xnor2_1 _06038_ (.A(_05166_),
    .B(_05167_),
    .Y(_05168_));
 sky130_fd_sc_hd__and3_1 _06039_ (.A(_05100_),
    .B(_05102_),
    .C(_05168_),
    .X(_05169_));
 sky130_fd_sc_hd__a21o_1 _06040_ (.A1(_05100_),
    .A2(_05102_),
    .B1(_05168_),
    .X(_05170_));
 sky130_fd_sc_hd__nand2b_1 _06041_ (.A_N(_05169_),
    .B(_05170_),
    .Y(_05171_));
 sky130_fd_sc_hd__xor2_1 _06042_ (.A(_05078_),
    .B(_05171_),
    .X(_05172_));
 sky130_fd_sc_hd__nand2_1 _06043_ (.A(_05096_),
    .B(_05098_),
    .Y(_05173_));
 sky130_fd_sc_hd__a21o_1 _06044_ (.A1(_05105_),
    .A2(_05112_),
    .B1(_05111_),
    .X(_05174_));
 sky130_fd_sc_hd__nand2_1 _06045_ (.A(net495),
    .B(net402),
    .Y(_05175_));
 sky130_fd_sc_hd__and4_1 _06046_ (.A(net480),
    .B(net492),
    .C(net417),
    .D(net409),
    .X(_05176_));
 sky130_fd_sc_hd__a22oi_1 _06047_ (.A1(net480),
    .A2(net417),
    .B1(net409),
    .B2(net492),
    .Y(_05177_));
 sky130_fd_sc_hd__nor2_1 _06048_ (.A(_05176_),
    .B(_05177_),
    .Y(_05178_));
 sky130_fd_sc_hd__xnor2_1 _06049_ (.A(_05175_),
    .B(_05178_),
    .Y(_05179_));
 sky130_fd_sc_hd__nand2_1 _06050_ (.A(net472),
    .B(net423),
    .Y(_05180_));
 sky130_fd_sc_hd__nand4_1 _06051_ (.A(net457),
    .B(net452),
    .C(net188),
    .D(net431),
    .Y(_05181_));
 sky130_fd_sc_hd__a22o_1 _06052_ (.A1(net452),
    .A2(net188),
    .B1(net431),
    .B2(net462),
    .X(_05182_));
 sky130_fd_sc_hd__nand3b_1 _06053_ (.A_N(_05180_),
    .B(_05181_),
    .C(_05182_),
    .Y(_05183_));
 sky130_fd_sc_hd__a21bo_1 _06054_ (.A1(_05181_),
    .A2(_05182_),
    .B1_N(_05180_),
    .X(_05184_));
 sky130_fd_sc_hd__a21bo_1 _06055_ (.A1(_05091_),
    .A2(_05092_),
    .B1_N(_05090_),
    .X(_05185_));
 sky130_fd_sc_hd__nand3_1 _06056_ (.A(_05183_),
    .B(_05184_),
    .C(_05185_),
    .Y(_05186_));
 sky130_fd_sc_hd__a21o_1 _06057_ (.A1(_05183_),
    .A2(_05184_),
    .B1(_05185_),
    .X(_05187_));
 sky130_fd_sc_hd__nand3_1 _06058_ (.A(_05179_),
    .B(_05186_),
    .C(_05187_),
    .Y(_05188_));
 sky130_fd_sc_hd__a21o_1 _06059_ (.A1(_05186_),
    .A2(_05187_),
    .B1(_05179_),
    .X(_05189_));
 sky130_fd_sc_hd__nand3_1 _06060_ (.A(_05174_),
    .B(_05188_),
    .C(_05189_),
    .Y(_05190_));
 sky130_fd_sc_hd__a21o_1 _06061_ (.A1(_05188_),
    .A2(_05189_),
    .B1(_05174_),
    .X(_05191_));
 sky130_fd_sc_hd__and3_1 _06062_ (.A(_05173_),
    .B(_05190_),
    .C(_05191_),
    .X(_05192_));
 sky130_fd_sc_hd__a21oi_1 _06063_ (.A1(_05190_),
    .A2(_05191_),
    .B1(_05173_),
    .Y(_05193_));
 sky130_fd_sc_hd__or2_1 _06064_ (.A(_05192_),
    .B(_05193_),
    .X(_05194_));
 sky130_fd_sc_hd__nand2_1 _06065_ (.A(_05107_),
    .B(_05110_),
    .Y(_05195_));
 sky130_fd_sc_hd__o21ba_1 _06066_ (.A1(_05116_),
    .A2(_05118_),
    .B1_N(_05115_),
    .X(_05196_));
 sky130_fd_sc_hd__nand2_1 _06067_ (.A(net195),
    .B(net446),
    .Y(_05197_));
 sky130_fd_sc_hd__and4_1 _06068_ (.A(net214),
    .B(net205),
    .C(net547),
    .D(net466),
    .X(_05198_));
 sky130_fd_sc_hd__a22oi_1 _06069_ (.A1(net205),
    .A2(net547),
    .B1(net466),
    .B2(net214),
    .Y(_05199_));
 sky130_fd_sc_hd__nor2_1 _06070_ (.A(_05198_),
    .B(_05199_),
    .Y(_05200_));
 sky130_fd_sc_hd__xnor2_1 _06071_ (.A(_05197_),
    .B(_05200_),
    .Y(_05201_));
 sky130_fd_sc_hd__nand2b_1 _06072_ (.A_N(_05196_),
    .B(_05201_),
    .Y(_05202_));
 sky130_fd_sc_hd__xnor2_1 _06073_ (.A(_05196_),
    .B(_05201_),
    .Y(_05203_));
 sky130_fd_sc_hd__nand2_1 _06074_ (.A(_05195_),
    .B(_05203_),
    .Y(_05204_));
 sky130_fd_sc_hd__xor2_1 _06075_ (.A(_05195_),
    .B(_05203_),
    .X(_05205_));
 sky130_fd_sc_hd__nand2_1 _06076_ (.A(net217),
    .B(net384),
    .Y(_05206_));
 sky130_fd_sc_hd__and4_1 _06077_ (.A(net241),
    .B(net232),
    .C(net302),
    .D(net226),
    .X(_05207_));
 sky130_fd_sc_hd__a22oi_1 _06078_ (.A1(net232),
    .A2(net302),
    .B1(net226),
    .B2(net241),
    .Y(_05208_));
 sky130_fd_sc_hd__nor2_1 _06079_ (.A(_05207_),
    .B(_05208_),
    .Y(_05209_));
 sky130_fd_sc_hd__xnor2_1 _06080_ (.A(_05206_),
    .B(_05209_),
    .Y(_05210_));
 sky130_fd_sc_hd__nand2_1 _06081_ (.A(net256),
    .B(net181),
    .Y(_05211_));
 sky130_fd_sc_hd__and4_1 _06082_ (.A(net439),
    .B(net345),
    .C(net171),
    .D(net163),
    .X(_05212_));
 sky130_fd_sc_hd__a22oi_2 _06083_ (.A1(net346),
    .A2(net171),
    .B1(net163),
    .B2(net439),
    .Y(_05213_));
 sky130_fd_sc_hd__or3_1 _06084_ (.A(_05211_),
    .B(_05212_),
    .C(_05213_),
    .X(_05214_));
 sky130_fd_sc_hd__o21ai_1 _06085_ (.A1(_05212_),
    .A2(_05213_),
    .B1(_05211_),
    .Y(_05215_));
 sky130_fd_sc_hd__o21bai_1 _06086_ (.A1(_05120_),
    .A2(_05122_),
    .B1_N(_05121_),
    .Y(_05216_));
 sky130_fd_sc_hd__nand3_1 _06087_ (.A(_05214_),
    .B(_05215_),
    .C(_05216_),
    .Y(_05217_));
 sky130_fd_sc_hd__a21o_1 _06088_ (.A1(_05214_),
    .A2(_05215_),
    .B1(_05216_),
    .X(_05218_));
 sky130_fd_sc_hd__nand3_1 _06089_ (.A(_05210_),
    .B(_05217_),
    .C(_05218_),
    .Y(_05219_));
 sky130_fd_sc_hd__a21o_1 _06090_ (.A1(_05217_),
    .A2(_05218_),
    .B1(_05210_),
    .X(_05220_));
 sky130_fd_sc_hd__a21bo_1 _06091_ (.A1(_05119_),
    .A2(_05127_),
    .B1_N(_05126_),
    .X(_05221_));
 sky130_fd_sc_hd__nand3_4 _06092_ (.A(_05219_),
    .B(_05220_),
    .C(_05221_),
    .Y(_05222_));
 sky130_fd_sc_hd__a21o_1 _06093_ (.A1(_05219_),
    .A2(_05220_),
    .B1(_05221_),
    .X(_05223_));
 sky130_fd_sc_hd__and3_1 _06094_ (.A(_05205_),
    .B(_05222_),
    .C(_05223_),
    .X(_05224_));
 sky130_fd_sc_hd__nand3_2 _06095_ (.A(_05205_),
    .B(_05222_),
    .C(_05223_),
    .Y(_05225_));
 sky130_fd_sc_hd__a21oi_1 _06096_ (.A1(_05222_),
    .A2(_05223_),
    .B1(_05205_),
    .Y(_05226_));
 sky130_fd_sc_hd__a211oi_2 _06097_ (.A1(_05131_),
    .A2(_05134_),
    .B1(_05224_),
    .C1(_05226_),
    .Y(_05227_));
 sky130_fd_sc_hd__o211a_1 _06098_ (.A1(_05224_),
    .A2(_05226_),
    .B1(_05131_),
    .C1(_05134_),
    .X(_05228_));
 sky130_fd_sc_hd__nor3_1 _06099_ (.A(_05194_),
    .B(_05227_),
    .C(_05228_),
    .Y(_05229_));
 sky130_fd_sc_hd__or3_1 _06100_ (.A(_05194_),
    .B(_05227_),
    .C(_05228_),
    .X(_05230_));
 sky130_fd_sc_hd__o21ai_1 _06101_ (.A1(_05227_),
    .A2(_05228_),
    .B1(_05194_),
    .Y(_05231_));
 sky130_fd_sc_hd__o211ai_2 _06102_ (.A1(_05136_),
    .A2(_05138_),
    .B1(_05230_),
    .C1(_05231_),
    .Y(_05232_));
 sky130_fd_sc_hd__a211o_1 _06103_ (.A1(_05230_),
    .A2(_05231_),
    .B1(_05136_),
    .C1(_05138_),
    .X(_05233_));
 sky130_fd_sc_hd__and3_1 _06104_ (.A(_05172_),
    .B(_05232_),
    .C(_05233_),
    .X(_05234_));
 sky130_fd_sc_hd__a21oi_1 _06105_ (.A1(_05232_),
    .A2(_05233_),
    .B1(_05172_),
    .Y(_05235_));
 sky130_fd_sc_hd__a211o_1 _06106_ (.A1(_05140_),
    .A2(_05142_),
    .B1(_05234_),
    .C1(_05235_),
    .X(_05236_));
 sky130_fd_sc_hd__inv_2 _06107_ (.A(_05236_),
    .Y(_05237_));
 sky130_fd_sc_hd__o211ai_1 _06108_ (.A1(_05234_),
    .A2(_05235_),
    .B1(_05140_),
    .C1(_05142_),
    .Y(_05238_));
 sky130_fd_sc_hd__and3_1 _06109_ (.A(_05081_),
    .B(_05236_),
    .C(_05238_),
    .X(_05239_));
 sky130_fd_sc_hd__a21oi_1 _06110_ (.A1(_05236_),
    .A2(_05238_),
    .B1(_05081_),
    .Y(_05240_));
 sky130_fd_sc_hd__a211o_1 _06111_ (.A1(_05144_),
    .A2(_05146_),
    .B1(_05239_),
    .C1(_05240_),
    .X(_05241_));
 sky130_fd_sc_hd__o211ai_1 _06112_ (.A1(_05239_),
    .A2(_05240_),
    .B1(_05144_),
    .C1(_05146_),
    .Y(_05242_));
 sky130_fd_sc_hd__and3_1 _06113_ (.A(_05148_),
    .B(_05241_),
    .C(_05242_),
    .X(_05243_));
 sky130_fd_sc_hd__a21oi_1 _06114_ (.A1(_05241_),
    .A2(_05242_),
    .B1(_05148_),
    .Y(_05244_));
 sky130_fd_sc_hd__nor2_1 _06115_ (.A(_05243_),
    .B(_05244_),
    .Y(_05245_));
 sky130_fd_sc_hd__or3_1 _06116_ (.A(_05153_),
    .B(_05243_),
    .C(_05244_),
    .X(_05246_));
 sky130_fd_sc_hd__xnor2_1 _06117_ (.A(_05153_),
    .B(_05245_),
    .Y(_05247_));
 sky130_fd_sc_hd__xnor2_1 _06118_ (.A(_05156_),
    .B(_05247_),
    .Y(net73));
 sky130_fd_sc_hd__nor2_1 _06119_ (.A(_05237_),
    .B(_05239_),
    .Y(_05248_));
 sky130_fd_sc_hd__o21a_1 _06120_ (.A1(_05078_),
    .A2(_05169_),
    .B1(_05170_),
    .X(_05249_));
 sky130_fd_sc_hd__and3b_1 _06121_ (.A_N(_05164_),
    .B(_05075_),
    .C(_05163_),
    .X(_05250_));
 sky130_fd_sc_hd__a31o_1 _06122_ (.A1(_05174_),
    .A2(_05188_),
    .A3(_05189_),
    .B1(_05192_),
    .X(_05251_));
 sky130_fd_sc_hd__or2_1 _06123_ (.A(_05158_),
    .B(_05160_),
    .X(_05252_));
 sky130_fd_sc_hd__o21ba_1 _06124_ (.A1(_05175_),
    .A2(_05177_),
    .B1_N(_05176_),
    .X(_05253_));
 sky130_fd_sc_hd__and4_1 _06125_ (.A(net499),
    .B(net519),
    .C(net394),
    .D(net378),
    .X(_05254_));
 sky130_fd_sc_hd__a22oi_1 _06126_ (.A1(net499),
    .A2(net394),
    .B1(net378),
    .B2(net519),
    .Y(_05255_));
 sky130_fd_sc_hd__nor2_1 _06127_ (.A(_05254_),
    .B(_05255_),
    .Y(_05256_));
 sky130_fd_sc_hd__nand2_1 _06128_ (.A(net604),
    .B(net370),
    .Y(_05257_));
 sky130_fd_sc_hd__xnor2_1 _06129_ (.A(_05256_),
    .B(_05257_),
    .Y(_05258_));
 sky130_fd_sc_hd__nand2b_1 _06130_ (.A_N(_05253_),
    .B(_05258_),
    .Y(_05259_));
 sky130_fd_sc_hd__xnor2_1 _06131_ (.A(_05253_),
    .B(_05258_),
    .Y(_05260_));
 sky130_fd_sc_hd__nand2_1 _06132_ (.A(_05252_),
    .B(_05260_),
    .Y(_05261_));
 sky130_fd_sc_hd__xnor2_1 _06133_ (.A(_05252_),
    .B(_05260_),
    .Y(_05262_));
 sky130_fd_sc_hd__o21ai_1 _06134_ (.A1(_05072_),
    .A2(_05164_),
    .B1(_05163_),
    .Y(_05263_));
 sky130_fd_sc_hd__xor2_1 _06135_ (.A(_05262_),
    .B(_05263_),
    .X(_05264_));
 sky130_fd_sc_hd__nand2_1 _06136_ (.A(net629),
    .B(net360),
    .Y(_05265_));
 sky130_fd_sc_hd__and3_1 _06137_ (.A(net629),
    .B(net360),
    .C(_05264_),
    .X(_05266_));
 sky130_fd_sc_hd__xor2_1 _06138_ (.A(_05264_),
    .B(_05265_),
    .X(_05267_));
 sky130_fd_sc_hd__and2b_1 _06139_ (.A_N(_05267_),
    .B(_05251_),
    .X(_05268_));
 sky130_fd_sc_hd__xnor2_1 _06140_ (.A(_05251_),
    .B(_05267_),
    .Y(_05269_));
 sky130_fd_sc_hd__xnor2_1 _06141_ (.A(_05250_),
    .B(_05269_),
    .Y(_05270_));
 sky130_fd_sc_hd__nand2_1 _06142_ (.A(_05186_),
    .B(_05188_),
    .Y(_05271_));
 sky130_fd_sc_hd__nand2_1 _06143_ (.A(net491),
    .B(net402),
    .Y(_05272_));
 sky130_fd_sc_hd__and4_1 _06144_ (.A(net483),
    .B(net475),
    .C(net417),
    .D(net409),
    .X(_05273_));
 sky130_fd_sc_hd__a22oi_1 _06145_ (.A1(net475),
    .A2(net418),
    .B1(net410),
    .B2(net483),
    .Y(_05274_));
 sky130_fd_sc_hd__nor2_1 _06146_ (.A(_05273_),
    .B(_05274_),
    .Y(_05275_));
 sky130_fd_sc_hd__xnor2_1 _06147_ (.A(_05272_),
    .B(_05275_),
    .Y(_05276_));
 sky130_fd_sc_hd__nand2_1 _06148_ (.A(net462),
    .B(net423),
    .Y(_05277_));
 sky130_fd_sc_hd__and4_1 _06149_ (.A(net452),
    .B(net446),
    .C(net188),
    .D(net431),
    .X(_05278_));
 sky130_fd_sc_hd__a22oi_1 _06150_ (.A1(net446),
    .A2(net188),
    .B1(net431),
    .B2(net455),
    .Y(_05279_));
 sky130_fd_sc_hd__nor2_1 _06151_ (.A(_05278_),
    .B(_05279_),
    .Y(_05280_));
 sky130_fd_sc_hd__xnor2_1 _06152_ (.A(_05277_),
    .B(_05280_),
    .Y(_05281_));
 sky130_fd_sc_hd__nand2_1 _06153_ (.A(_05181_),
    .B(_05183_),
    .Y(_05282_));
 sky130_fd_sc_hd__and2_1 _06154_ (.A(_05281_),
    .B(_05282_),
    .X(_05283_));
 sky130_fd_sc_hd__xor2_1 _06155_ (.A(_05281_),
    .B(_05282_),
    .X(_05284_));
 sky130_fd_sc_hd__and2_1 _06156_ (.A(_05276_),
    .B(_05284_),
    .X(_05285_));
 sky130_fd_sc_hd__xnor2_1 _06157_ (.A(_05276_),
    .B(_05284_),
    .Y(_05286_));
 sky130_fd_sc_hd__a21o_1 _06158_ (.A1(_05202_),
    .A2(_05204_),
    .B1(_05286_),
    .X(_05287_));
 sky130_fd_sc_hd__nand3_1 _06159_ (.A(_05202_),
    .B(_05204_),
    .C(_05286_),
    .Y(_05288_));
 sky130_fd_sc_hd__and3_1 _06160_ (.A(_05271_),
    .B(_05287_),
    .C(_05288_),
    .X(_05289_));
 sky130_fd_sc_hd__nand3_1 _06161_ (.A(_05271_),
    .B(_05287_),
    .C(_05288_),
    .Y(_05290_));
 sky130_fd_sc_hd__a21oi_1 _06162_ (.A1(_05287_),
    .A2(_05288_),
    .B1(_05271_),
    .Y(_05291_));
 sky130_fd_sc_hd__o21ba_1 _06163_ (.A1(_05197_),
    .A2(_05199_),
    .B1_N(_05198_),
    .X(_05292_));
 sky130_fd_sc_hd__o21ba_1 _06164_ (.A1(_05206_),
    .A2(_05208_),
    .B1_N(_05207_),
    .X(_05293_));
 sky130_fd_sc_hd__nand2_1 _06165_ (.A(net195),
    .B(net547),
    .Y(_05294_));
 sky130_fd_sc_hd__and4_1 _06166_ (.A(net212),
    .B(net203),
    .C(net466),
    .D(net385),
    .X(_05295_));
 sky130_fd_sc_hd__a22oi_1 _06167_ (.A1(net203),
    .A2(net466),
    .B1(net385),
    .B2(net212),
    .Y(_05296_));
 sky130_fd_sc_hd__nor2_1 _06168_ (.A(_05295_),
    .B(_05296_),
    .Y(_05297_));
 sky130_fd_sc_hd__xnor2_1 _06169_ (.A(_05294_),
    .B(_05297_),
    .Y(_05298_));
 sky130_fd_sc_hd__nand2b_1 _06170_ (.A_N(_05293_),
    .B(_05298_),
    .Y(_05299_));
 sky130_fd_sc_hd__xnor2_1 _06171_ (.A(_05293_),
    .B(_05298_),
    .Y(_05300_));
 sky130_fd_sc_hd__nand2b_1 _06172_ (.A_N(_05292_),
    .B(_05300_),
    .Y(_05301_));
 sky130_fd_sc_hd__xnor2_1 _06173_ (.A(_05292_),
    .B(_05300_),
    .Y(_05302_));
 sky130_fd_sc_hd__nand2_1 _06174_ (.A(net217),
    .B(net302),
    .Y(_05303_));
 sky130_fd_sc_hd__and4_1 _06175_ (.A(net240),
    .B(net233),
    .C(net226),
    .D(net179),
    .X(_05304_));
 sky130_fd_sc_hd__a22oi_1 _06176_ (.A1(net232),
    .A2(net226),
    .B1(net179),
    .B2(net240),
    .Y(_05305_));
 sky130_fd_sc_hd__nor2_1 _06177_ (.A(_05304_),
    .B(_05305_),
    .Y(_05306_));
 sky130_fd_sc_hd__xnor2_1 _06178_ (.A(_05303_),
    .B(_05306_),
    .Y(_00000_));
 sky130_fd_sc_hd__nand2_1 _06179_ (.A(net256),
    .B(net171),
    .Y(_00001_));
 sky130_fd_sc_hd__and4_1 _06180_ (.A(net437),
    .B(net345),
    .C(net163),
    .D(net622),
    .X(_00002_));
 sky130_fd_sc_hd__a22oi_2 _06181_ (.A1(net345),
    .A2(net163),
    .B1(net622),
    .B2(net437),
    .Y(_00003_));
 sky130_fd_sc_hd__or3_1 _06182_ (.A(_00001_),
    .B(_00002_),
    .C(_00003_),
    .X(_00004_));
 sky130_fd_sc_hd__o21ai_1 _06183_ (.A1(_00002_),
    .A2(_00003_),
    .B1(_00001_),
    .Y(_00005_));
 sky130_fd_sc_hd__o21bai_1 _06184_ (.A1(_05211_),
    .A2(_05213_),
    .B1_N(_05212_),
    .Y(_00006_));
 sky130_fd_sc_hd__nand3_1 _06185_ (.A(_00004_),
    .B(_00005_),
    .C(_00006_),
    .Y(_00007_));
 sky130_fd_sc_hd__a21o_1 _06186_ (.A1(_00004_),
    .A2(_00005_),
    .B1(_00006_),
    .X(_00008_));
 sky130_fd_sc_hd__nand3_1 _06187_ (.A(_00000_),
    .B(_00007_),
    .C(_00008_),
    .Y(_00009_));
 sky130_fd_sc_hd__a21o_1 _06188_ (.A1(_00007_),
    .A2(_00008_),
    .B1(_00000_),
    .X(_00010_));
 sky130_fd_sc_hd__a21bo_1 _06189_ (.A1(_05210_),
    .A2(_05218_),
    .B1_N(_05217_),
    .X(_00011_));
 sky130_fd_sc_hd__nand3_4 _06190_ (.A(_00009_),
    .B(_00010_),
    .C(_00011_),
    .Y(_00012_));
 sky130_fd_sc_hd__a21o_1 _06191_ (.A1(_00009_),
    .A2(_00010_),
    .B1(_00011_),
    .X(_00013_));
 sky130_fd_sc_hd__and3_1 _06192_ (.A(_05302_),
    .B(_00012_),
    .C(_00013_),
    .X(_00014_));
 sky130_fd_sc_hd__nand3_2 _06193_ (.A(_05302_),
    .B(_00012_),
    .C(_00013_),
    .Y(_00015_));
 sky130_fd_sc_hd__a21oi_2 _06194_ (.A1(_00012_),
    .A2(_00013_),
    .B1(_05302_),
    .Y(_00016_));
 sky130_fd_sc_hd__a211oi_4 _06195_ (.A1(_05222_),
    .A2(_05225_),
    .B1(_00014_),
    .C1(_00016_),
    .Y(_00017_));
 sky130_fd_sc_hd__o211a_1 _06196_ (.A1(_00014_),
    .A2(_00016_),
    .B1(_05222_),
    .C1(_05225_),
    .X(_00018_));
 sky130_fd_sc_hd__nor4_1 _06197_ (.A(_05289_),
    .B(_05291_),
    .C(_00017_),
    .D(_00018_),
    .Y(_00019_));
 sky130_fd_sc_hd__or4_1 _06198_ (.A(_05289_),
    .B(_05291_),
    .C(_00017_),
    .D(_00018_),
    .X(_00020_));
 sky130_fd_sc_hd__o22ai_1 _06199_ (.A1(_05289_),
    .A2(_05291_),
    .B1(_00017_),
    .B2(_00018_),
    .Y(_00021_));
 sky130_fd_sc_hd__o211a_1 _06200_ (.A1(_05227_),
    .A2(_05229_),
    .B1(_00020_),
    .C1(_00021_),
    .X(_00022_));
 sky130_fd_sc_hd__a211oi_1 _06201_ (.A1(_00020_),
    .A2(_00021_),
    .B1(_05227_),
    .C1(_05229_),
    .Y(_00023_));
 sky130_fd_sc_hd__or3_1 _06202_ (.A(_05270_),
    .B(_00022_),
    .C(_00023_),
    .X(_00024_));
 sky130_fd_sc_hd__o21ai_1 _06203_ (.A1(_00022_),
    .A2(_00023_),
    .B1(_05270_),
    .Y(_00025_));
 sky130_fd_sc_hd__a21bo_1 _06204_ (.A1(_05172_),
    .A2(_05233_),
    .B1_N(_05232_),
    .X(_00026_));
 sky130_fd_sc_hd__and3_1 _06205_ (.A(_00024_),
    .B(_00025_),
    .C(_00026_),
    .X(_00027_));
 sky130_fd_sc_hd__a21oi_1 _06206_ (.A1(_00024_),
    .A2(_00025_),
    .B1(_00026_),
    .Y(_00028_));
 sky130_fd_sc_hd__nor3_1 _06207_ (.A(_05249_),
    .B(_00027_),
    .C(_00028_),
    .Y(_00029_));
 sky130_fd_sc_hd__o21a_1 _06208_ (.A1(_00027_),
    .A2(_00028_),
    .B1(_05249_),
    .X(_00030_));
 sky130_fd_sc_hd__nor2_1 _06209_ (.A(_00029_),
    .B(_00030_),
    .Y(_00031_));
 sky130_fd_sc_hd__and2b_1 _06210_ (.A_N(_05248_),
    .B(_00031_),
    .X(_00032_));
 sky130_fd_sc_hd__xnor2_1 _06211_ (.A(_05248_),
    .B(_00031_),
    .Y(_00033_));
 sky130_fd_sc_hd__and2b_1 _06212_ (.A_N(_05241_),
    .B(_00033_),
    .X(_00034_));
 sky130_fd_sc_hd__xnor2_1 _06213_ (.A(_05241_),
    .B(_00033_),
    .Y(_00035_));
 sky130_fd_sc_hd__and2_1 _06214_ (.A(_05243_),
    .B(_00035_),
    .X(_00036_));
 sky130_fd_sc_hd__nor2_1 _06215_ (.A(_05243_),
    .B(_00035_),
    .Y(_00037_));
 sky130_fd_sc_hd__nor2_1 _06216_ (.A(_00036_),
    .B(_00037_),
    .Y(_00038_));
 sky130_fd_sc_hd__o21ai_1 _06217_ (.A1(_05066_),
    .A2(_05245_),
    .B1(_05150_),
    .Y(_00039_));
 sky130_fd_sc_hd__o21ai_1 _06218_ (.A1(_05071_),
    .A2(_00039_),
    .B1(_05246_),
    .Y(_00040_));
 sky130_fd_sc_hd__and2_1 _06219_ (.A(_05154_),
    .B(_05245_),
    .X(_00041_));
 sky130_fd_sc_hd__inv_2 _06220_ (.A(_00041_),
    .Y(_00042_));
 sky130_fd_sc_hd__o21ba_1 _06221_ (.A1(_05070_),
    .A2(_00042_),
    .B1_N(_00040_),
    .X(_00043_));
 sky130_fd_sc_hd__and2b_1 _06222_ (.A_N(_00043_),
    .B(_00038_),
    .X(_00044_));
 sky130_fd_sc_hd__xnor2_1 _06223_ (.A(_00038_),
    .B(_00043_),
    .Y(net74));
 sky130_fd_sc_hd__a21o_1 _06224_ (.A1(_05250_),
    .A2(_05269_),
    .B1(_05268_),
    .X(_00045_));
 sky130_fd_sc_hd__o21ba_1 _06225_ (.A1(_05262_),
    .A2(_05263_),
    .B1_N(_05266_),
    .X(_00046_));
 sky130_fd_sc_hd__a22o_1 _06226_ (.A1(net604),
    .A2(net360),
    .B1(net352),
    .B2(net629),
    .X(_00047_));
 sky130_fd_sc_hd__nand2_1 _06227_ (.A(net604),
    .B(net356),
    .Y(_00048_));
 sky130_fd_sc_hd__nor2_1 _06228_ (.A(_05265_),
    .B(_00048_),
    .Y(_00049_));
 sky130_fd_sc_hd__or2_1 _06229_ (.A(_05265_),
    .B(_00048_),
    .X(_00050_));
 sky130_fd_sc_hd__a31o_1 _06230_ (.A1(net604),
    .A2(net370),
    .A3(_05256_),
    .B1(_05254_),
    .X(_00051_));
 sky130_fd_sc_hd__o21ba_1 _06231_ (.A1(_05272_),
    .A2(_05274_),
    .B1_N(_05273_),
    .X(_00052_));
 sky130_fd_sc_hd__and4_1 _06232_ (.A(net491),
    .B(net499),
    .C(net394),
    .D(net378),
    .X(_00053_));
 sky130_fd_sc_hd__a22oi_1 _06233_ (.A1(net491),
    .A2(net395),
    .B1(net378),
    .B2(net499),
    .Y(_00054_));
 sky130_fd_sc_hd__nor2_1 _06234_ (.A(_00053_),
    .B(_00054_),
    .Y(_00055_));
 sky130_fd_sc_hd__nand2_1 _06235_ (.A(net519),
    .B(net370),
    .Y(_00056_));
 sky130_fd_sc_hd__xnor2_1 _06236_ (.A(_00055_),
    .B(_00056_),
    .Y(_00057_));
 sky130_fd_sc_hd__nand2b_1 _06237_ (.A_N(_00052_),
    .B(_00057_),
    .Y(_00058_));
 sky130_fd_sc_hd__xnor2_1 _06238_ (.A(_00052_),
    .B(_00057_),
    .Y(_00059_));
 sky130_fd_sc_hd__nand2_1 _06239_ (.A(_00051_),
    .B(_00059_),
    .Y(_00060_));
 sky130_fd_sc_hd__xnor2_1 _06240_ (.A(_00051_),
    .B(_00059_),
    .Y(_00061_));
 sky130_fd_sc_hd__a21o_1 _06241_ (.A1(_05259_),
    .A2(_05261_),
    .B1(_00061_),
    .X(_00062_));
 sky130_fd_sc_hd__nand3_1 _06242_ (.A(_05259_),
    .B(_05261_),
    .C(_00061_),
    .Y(_00063_));
 sky130_fd_sc_hd__and4_1 _06243_ (.A(_00047_),
    .B(_00050_),
    .C(_00062_),
    .D(_00063_),
    .X(_00064_));
 sky130_fd_sc_hd__nand4_1 _06244_ (.A(_00047_),
    .B(_00050_),
    .C(_00062_),
    .D(_00063_),
    .Y(_00065_));
 sky130_fd_sc_hd__a22oi_1 _06245_ (.A1(_00047_),
    .A2(_00050_),
    .B1(_00062_),
    .B2(_00063_),
    .Y(_00066_));
 sky130_fd_sc_hd__a211oi_1 _06246_ (.A1(_05287_),
    .A2(_05290_),
    .B1(_00064_),
    .C1(_00066_),
    .Y(_00067_));
 sky130_fd_sc_hd__o211a_1 _06247_ (.A1(_00064_),
    .A2(_00066_),
    .B1(_05287_),
    .C1(_05290_),
    .X(_00068_));
 sky130_fd_sc_hd__nor3_1 _06248_ (.A(_00046_),
    .B(_00067_),
    .C(_00068_),
    .Y(_00069_));
 sky130_fd_sc_hd__o21a_1 _06249_ (.A1(_00067_),
    .A2(_00068_),
    .B1(_00046_),
    .X(_00070_));
 sky130_fd_sc_hd__nand2_1 _06250_ (.A(net483),
    .B(net402),
    .Y(_00071_));
 sky130_fd_sc_hd__and4_1 _06251_ (.A(net475),
    .B(net460),
    .C(net418),
    .D(net410),
    .X(_00072_));
 sky130_fd_sc_hd__a22oi_1 _06252_ (.A1(net460),
    .A2(net418),
    .B1(net410),
    .B2(net475),
    .Y(_00073_));
 sky130_fd_sc_hd__nor2_1 _06253_ (.A(_00072_),
    .B(_00073_),
    .Y(_00074_));
 sky130_fd_sc_hd__xnor2_1 _06254_ (.A(_00071_),
    .B(_00074_),
    .Y(_00075_));
 sky130_fd_sc_hd__nand2_1 _06255_ (.A(net453),
    .B(net423),
    .Y(_00076_));
 sky130_fd_sc_hd__and4_1 _06256_ (.A(net548),
    .B(net447),
    .C(net188),
    .D(net431),
    .X(_00077_));
 sky130_fd_sc_hd__a22oi_1 _06257_ (.A1(net548),
    .A2(net188),
    .B1(net431),
    .B2(net447),
    .Y(_00078_));
 sky130_fd_sc_hd__nor2_1 _06258_ (.A(_00077_),
    .B(_00078_),
    .Y(_00079_));
 sky130_fd_sc_hd__xnor2_1 _06259_ (.A(_00076_),
    .B(_00079_),
    .Y(_00080_));
 sky130_fd_sc_hd__o21ba_1 _06260_ (.A1(_05277_),
    .A2(_05279_),
    .B1_N(_05278_),
    .X(_00081_));
 sky130_fd_sc_hd__and2b_1 _06261_ (.A_N(_00081_),
    .B(_00080_),
    .X(_00082_));
 sky130_fd_sc_hd__xnor2_1 _06262_ (.A(_00080_),
    .B(_00081_),
    .Y(_00083_));
 sky130_fd_sc_hd__and2_1 _06263_ (.A(_00075_),
    .B(_00083_),
    .X(_00084_));
 sky130_fd_sc_hd__xnor2_1 _06264_ (.A(_00075_),
    .B(_00083_),
    .Y(_00085_));
 sky130_fd_sc_hd__a21o_2 _06265_ (.A1(_05299_),
    .A2(_05301_),
    .B1(_00085_),
    .X(_00086_));
 sky130_fd_sc_hd__nand3_1 _06266_ (.A(_05299_),
    .B(_05301_),
    .C(_00085_),
    .Y(_00087_));
 sky130_fd_sc_hd__o211a_1 _06267_ (.A1(_05283_),
    .A2(_05285_),
    .B1(_00086_),
    .C1(_00087_),
    .X(_00088_));
 sky130_fd_sc_hd__o211ai_2 _06268_ (.A1(_05283_),
    .A2(_05285_),
    .B1(_00086_),
    .C1(_00087_),
    .Y(_00089_));
 sky130_fd_sc_hd__a211oi_2 _06269_ (.A1(_00086_),
    .A2(_00087_),
    .B1(_05283_),
    .C1(_05285_),
    .Y(_00090_));
 sky130_fd_sc_hd__o21ba_1 _06270_ (.A1(_05294_),
    .A2(_05296_),
    .B1_N(_05295_),
    .X(_00091_));
 sky130_fd_sc_hd__o21ba_1 _06271_ (.A1(_05303_),
    .A2(_05305_),
    .B1_N(_05304_),
    .X(_00092_));
 sky130_fd_sc_hd__nand2_1 _06272_ (.A(net195),
    .B(net466),
    .Y(_00093_));
 sky130_fd_sc_hd__and4_1 _06273_ (.A(net212),
    .B(net203),
    .C(net385),
    .D(net300),
    .X(_00094_));
 sky130_fd_sc_hd__a22oi_1 _06274_ (.A1(net203),
    .A2(net385),
    .B1(net300),
    .B2(net212),
    .Y(_00095_));
 sky130_fd_sc_hd__nor2_1 _06275_ (.A(_00094_),
    .B(_00095_),
    .Y(_00096_));
 sky130_fd_sc_hd__xnor2_1 _06276_ (.A(_00093_),
    .B(_00096_),
    .Y(_00097_));
 sky130_fd_sc_hd__nand2b_1 _06277_ (.A_N(_00092_),
    .B(_00097_),
    .Y(_00098_));
 sky130_fd_sc_hd__xnor2_1 _06278_ (.A(_00092_),
    .B(_00097_),
    .Y(_00099_));
 sky130_fd_sc_hd__nand2b_1 _06279_ (.A_N(_00091_),
    .B(_00099_),
    .Y(_00100_));
 sky130_fd_sc_hd__xnor2_1 _06280_ (.A(_00091_),
    .B(_00099_),
    .Y(_00101_));
 sky130_fd_sc_hd__nand2_1 _06281_ (.A(net217),
    .B(net226),
    .Y(_00102_));
 sky130_fd_sc_hd__and4_1 _06282_ (.A(net241),
    .B(net232),
    .C(net179),
    .D(net171),
    .X(_00103_));
 sky130_fd_sc_hd__a22oi_1 _06283_ (.A1(net232),
    .A2(net179),
    .B1(net171),
    .B2(net241),
    .Y(_00104_));
 sky130_fd_sc_hd__nor2_1 _06284_ (.A(_00103_),
    .B(_00104_),
    .Y(_00105_));
 sky130_fd_sc_hd__xnor2_1 _06285_ (.A(_00102_),
    .B(_00105_),
    .Y(_00106_));
 sky130_fd_sc_hd__nand2_1 _06286_ (.A(net256),
    .B(net163),
    .Y(_00107_));
 sky130_fd_sc_hd__and4_1 _06287_ (.A(net437),
    .B(net345),
    .C(net622),
    .D(net614),
    .X(_00108_));
 sky130_fd_sc_hd__a22oi_2 _06288_ (.A1(net345),
    .A2(net622),
    .B1(net614),
    .B2(net437),
    .Y(_00109_));
 sky130_fd_sc_hd__or3_1 _06289_ (.A(_00107_),
    .B(_00108_),
    .C(_00109_),
    .X(_00110_));
 sky130_fd_sc_hd__o21ai_1 _06290_ (.A1(_00108_),
    .A2(_00109_),
    .B1(_00107_),
    .Y(_00111_));
 sky130_fd_sc_hd__o21bai_1 _06291_ (.A1(_00001_),
    .A2(_00003_),
    .B1_N(_00002_),
    .Y(_00112_));
 sky130_fd_sc_hd__nand3_1 _06292_ (.A(_00110_),
    .B(_00111_),
    .C(_00112_),
    .Y(_00113_));
 sky130_fd_sc_hd__a21o_1 _06293_ (.A1(_00110_),
    .A2(_00111_),
    .B1(_00112_),
    .X(_00114_));
 sky130_fd_sc_hd__nand3_1 _06294_ (.A(_00106_),
    .B(_00113_),
    .C(_00114_),
    .Y(_00115_));
 sky130_fd_sc_hd__a21o_1 _06295_ (.A1(_00113_),
    .A2(_00114_),
    .B1(_00106_),
    .X(_00116_));
 sky130_fd_sc_hd__a21bo_1 _06296_ (.A1(_00000_),
    .A2(_00008_),
    .B1_N(_00007_),
    .X(_00117_));
 sky130_fd_sc_hd__nand3_4 _06297_ (.A(_00115_),
    .B(_00116_),
    .C(_00117_),
    .Y(_00118_));
 sky130_fd_sc_hd__a21o_1 _06298_ (.A1(_00115_),
    .A2(_00116_),
    .B1(_00117_),
    .X(_00119_));
 sky130_fd_sc_hd__and3_1 _06299_ (.A(_00101_),
    .B(_00118_),
    .C(_00119_),
    .X(_00120_));
 sky130_fd_sc_hd__nand3_2 _06300_ (.A(_00101_),
    .B(_00118_),
    .C(_00119_),
    .Y(_00121_));
 sky130_fd_sc_hd__a21oi_2 _06301_ (.A1(_00118_),
    .A2(_00119_),
    .B1(_00101_),
    .Y(_00122_));
 sky130_fd_sc_hd__a211oi_4 _06302_ (.A1(_00012_),
    .A2(_00015_),
    .B1(_00120_),
    .C1(_00122_),
    .Y(_00123_));
 sky130_fd_sc_hd__o211a_1 _06303_ (.A1(_00120_),
    .A2(_00122_),
    .B1(_00012_),
    .C1(_00015_),
    .X(_00124_));
 sky130_fd_sc_hd__nor4_1 _06304_ (.A(_00088_),
    .B(_00090_),
    .C(_00123_),
    .D(_00124_),
    .Y(_00125_));
 sky130_fd_sc_hd__or4_1 _06305_ (.A(_00088_),
    .B(_00090_),
    .C(_00123_),
    .D(_00124_),
    .X(_00126_));
 sky130_fd_sc_hd__o22ai_2 _06306_ (.A1(_00088_),
    .A2(_00090_),
    .B1(_00123_),
    .B2(_00124_),
    .Y(_00127_));
 sky130_fd_sc_hd__o211ai_2 _06307_ (.A1(_00017_),
    .A2(net151),
    .B1(_00126_),
    .C1(_00127_),
    .Y(_00128_));
 sky130_fd_sc_hd__a211o_1 _06308_ (.A1(_00126_),
    .A2(_00127_),
    .B1(_00017_),
    .C1(_00019_),
    .X(_00129_));
 sky130_fd_sc_hd__or4bb_2 _06309_ (.A(_00069_),
    .B(_00070_),
    .C_N(_00128_),
    .D_N(_00129_),
    .X(_00130_));
 sky130_fd_sc_hd__a2bb2o_1 _06310_ (.A1_N(_00069_),
    .A2_N(_00070_),
    .B1(_00128_),
    .B2(_00129_),
    .X(_00131_));
 sky130_fd_sc_hd__nand2_1 _06311_ (.A(_00130_),
    .B(_00131_),
    .Y(_00132_));
 sky130_fd_sc_hd__nand2b_1 _06312_ (.A_N(_00022_),
    .B(_00024_),
    .Y(_00133_));
 sky130_fd_sc_hd__xnor2_1 _06313_ (.A(_00132_),
    .B(_00133_),
    .Y(_00134_));
 sky130_fd_sc_hd__xnor2_1 _06314_ (.A(_00045_),
    .B(_00134_),
    .Y(_00135_));
 sky130_fd_sc_hd__nor2_1 _06315_ (.A(_00027_),
    .B(_00029_),
    .Y(_00136_));
 sky130_fd_sc_hd__or2_1 _06316_ (.A(_00135_),
    .B(_00136_),
    .X(_00137_));
 sky130_fd_sc_hd__xor2_1 _06317_ (.A(_00135_),
    .B(_00136_),
    .X(_00138_));
 sky130_fd_sc_hd__and2_1 _06318_ (.A(_00032_),
    .B(_00138_),
    .X(_00139_));
 sky130_fd_sc_hd__nor2_1 _06319_ (.A(_00032_),
    .B(_00138_),
    .Y(_00140_));
 sky130_fd_sc_hd__nor2_1 _06320_ (.A(_00139_),
    .B(_00140_),
    .Y(_00141_));
 sky130_fd_sc_hd__xor2_1 _06321_ (.A(_00034_),
    .B(_00141_),
    .X(_00142_));
 sky130_fd_sc_hd__nor2_1 _06322_ (.A(_00036_),
    .B(_00044_),
    .Y(_00143_));
 sky130_fd_sc_hd__xnor2_1 _06323_ (.A(_00142_),
    .B(_00143_),
    .Y(net75));
 sky130_fd_sc_hd__nor2_1 _06324_ (.A(_00067_),
    .B(_00069_),
    .Y(_00144_));
 sky130_fd_sc_hd__and4_1 _06325_ (.A(net519),
    .B(net604),
    .C(net364),
    .D(net356),
    .X(_00145_));
 sky130_fd_sc_hd__nand2_1 _06326_ (.A(net519),
    .B(net364),
    .Y(_00146_));
 sky130_fd_sc_hd__a21oi_1 _06327_ (.A1(_00048_),
    .A2(_00146_),
    .B1(_00145_),
    .Y(_00147_));
 sky130_fd_sc_hd__nand2_1 _06328_ (.A(net629),
    .B(net338),
    .Y(_00148_));
 sky130_fd_sc_hd__xnor2_1 _06329_ (.A(_00147_),
    .B(_00148_),
    .Y(_00149_));
 sky130_fd_sc_hd__and2_1 _06330_ (.A(_00049_),
    .B(_00149_),
    .X(_00150_));
 sky130_fd_sc_hd__nor2_1 _06331_ (.A(_00049_),
    .B(_00149_),
    .Y(_00151_));
 sky130_fd_sc_hd__or2_1 _06332_ (.A(_00150_),
    .B(_00151_),
    .X(_00152_));
 sky130_fd_sc_hd__a31o_1 _06333_ (.A1(net519),
    .A2(net370),
    .A3(_00055_),
    .B1(_00053_),
    .X(_00153_));
 sky130_fd_sc_hd__o21ba_1 _06334_ (.A1(_00071_),
    .A2(_00073_),
    .B1_N(_00072_),
    .X(_00154_));
 sky130_fd_sc_hd__and4_1 _06335_ (.A(net483),
    .B(net491),
    .C(net395),
    .D(net379),
    .X(_00155_));
 sky130_fd_sc_hd__a22oi_1 _06336_ (.A1(net483),
    .A2(net395),
    .B1(net379),
    .B2(net491),
    .Y(_00156_));
 sky130_fd_sc_hd__nor2_1 _06337_ (.A(_00155_),
    .B(_00156_),
    .Y(_00157_));
 sky130_fd_sc_hd__nand2_1 _06338_ (.A(net499),
    .B(net370),
    .Y(_00158_));
 sky130_fd_sc_hd__xnor2_1 _06339_ (.A(_00157_),
    .B(_00158_),
    .Y(_00159_));
 sky130_fd_sc_hd__nand2b_1 _06340_ (.A_N(_00154_),
    .B(_00159_),
    .Y(_00160_));
 sky130_fd_sc_hd__xnor2_1 _06341_ (.A(_00154_),
    .B(_00159_),
    .Y(_00161_));
 sky130_fd_sc_hd__nand2_1 _06342_ (.A(_00153_),
    .B(_00161_),
    .Y(_00162_));
 sky130_fd_sc_hd__xnor2_1 _06343_ (.A(_00153_),
    .B(_00161_),
    .Y(_00163_));
 sky130_fd_sc_hd__a21oi_2 _06344_ (.A1(_00058_),
    .A2(_00060_),
    .B1(_00163_),
    .Y(_00164_));
 sky130_fd_sc_hd__inv_2 _06345_ (.A(_00164_),
    .Y(_00165_));
 sky130_fd_sc_hd__and3_1 _06346_ (.A(_00058_),
    .B(_00060_),
    .C(_00163_),
    .X(_00166_));
 sky130_fd_sc_hd__nor3_1 _06347_ (.A(_00152_),
    .B(_00164_),
    .C(_00166_),
    .Y(_00167_));
 sky130_fd_sc_hd__or3_1 _06348_ (.A(_00152_),
    .B(_00164_),
    .C(_00166_),
    .X(_00168_));
 sky130_fd_sc_hd__o21a_1 _06349_ (.A1(_00164_),
    .A2(_00166_),
    .B1(_00152_),
    .X(_00169_));
 sky130_fd_sc_hd__a211oi_2 _06350_ (.A1(_00086_),
    .A2(_00089_),
    .B1(_00167_),
    .C1(_00169_),
    .Y(_00170_));
 sky130_fd_sc_hd__o211a_1 _06351_ (.A1(_00167_),
    .A2(_00169_),
    .B1(_00086_),
    .C1(_00089_),
    .X(_00171_));
 sky130_fd_sc_hd__a211oi_2 _06352_ (.A1(_00062_),
    .A2(_00065_),
    .B1(_00170_),
    .C1(_00171_),
    .Y(_00172_));
 sky130_fd_sc_hd__o211a_1 _06353_ (.A1(_00170_),
    .A2(_00171_),
    .B1(_00062_),
    .C1(_00065_),
    .X(_00173_));
 sky130_fd_sc_hd__nand2_1 _06354_ (.A(net475),
    .B(net402),
    .Y(_00174_));
 sky130_fd_sc_hd__and4_1 _06355_ (.A(net460),
    .B(net453),
    .C(net418),
    .D(net410),
    .X(_00175_));
 sky130_fd_sc_hd__a22oi_1 _06356_ (.A1(net453),
    .A2(net418),
    .B1(net410),
    .B2(net460),
    .Y(_00176_));
 sky130_fd_sc_hd__nor2_1 _06357_ (.A(_00175_),
    .B(_00176_),
    .Y(_00177_));
 sky130_fd_sc_hd__xnor2_1 _06358_ (.A(_00174_),
    .B(_00177_),
    .Y(_00178_));
 sky130_fd_sc_hd__nand2_1 _06359_ (.A(net447),
    .B(net424),
    .Y(_00179_));
 sky130_fd_sc_hd__and4_1 _06360_ (.A(net548),
    .B(net189),
    .C(net431),
    .D(net467),
    .X(_00180_));
 sky130_fd_sc_hd__a22oi_1 _06361_ (.A1(net548),
    .A2(net431),
    .B1(net467),
    .B2(net189),
    .Y(_00181_));
 sky130_fd_sc_hd__nor2_1 _06362_ (.A(_00180_),
    .B(_00181_),
    .Y(_00182_));
 sky130_fd_sc_hd__xnor2_1 _06363_ (.A(_00179_),
    .B(_00182_),
    .Y(_00183_));
 sky130_fd_sc_hd__o21ba_1 _06364_ (.A1(_00076_),
    .A2(_00078_),
    .B1_N(_00077_),
    .X(_00184_));
 sky130_fd_sc_hd__and2b_1 _06365_ (.A_N(_00184_),
    .B(_00183_),
    .X(_00185_));
 sky130_fd_sc_hd__xnor2_1 _06366_ (.A(_00183_),
    .B(_00184_),
    .Y(_00186_));
 sky130_fd_sc_hd__and2_1 _06367_ (.A(_00178_),
    .B(_00186_),
    .X(_00187_));
 sky130_fd_sc_hd__xnor2_1 _06368_ (.A(_00178_),
    .B(_00186_),
    .Y(_00188_));
 sky130_fd_sc_hd__a21o_2 _06369_ (.A1(_00098_),
    .A2(_00100_),
    .B1(_00188_),
    .X(_00189_));
 sky130_fd_sc_hd__nand3_2 _06370_ (.A(_00098_),
    .B(_00100_),
    .C(_00188_),
    .Y(_00190_));
 sky130_fd_sc_hd__o211a_1 _06371_ (.A1(_00082_),
    .A2(_00084_),
    .B1(_00189_),
    .C1(_00190_),
    .X(_00191_));
 sky130_fd_sc_hd__o211ai_2 _06372_ (.A1(_00082_),
    .A2(_00084_),
    .B1(_00189_),
    .C1(_00190_),
    .Y(_00192_));
 sky130_fd_sc_hd__a211oi_2 _06373_ (.A1(_00189_),
    .A2(_00190_),
    .B1(_00082_),
    .C1(_00084_),
    .Y(_00193_));
 sky130_fd_sc_hd__o21ba_1 _06374_ (.A1(_00093_),
    .A2(_00095_),
    .B1_N(_00094_),
    .X(_00194_));
 sky130_fd_sc_hd__o21ba_1 _06375_ (.A1(_00102_),
    .A2(_00104_),
    .B1_N(_00103_),
    .X(_00195_));
 sky130_fd_sc_hd__and4_1 _06376_ (.A(net212),
    .B(net204),
    .C(net300),
    .D(net224),
    .X(_00196_));
 sky130_fd_sc_hd__a22oi_1 _06377_ (.A1(net204),
    .A2(net300),
    .B1(net224),
    .B2(net213),
    .Y(_00197_));
 sky130_fd_sc_hd__nor2_1 _06378_ (.A(_00196_),
    .B(_00197_),
    .Y(_00198_));
 sky130_fd_sc_hd__nand2_1 _06379_ (.A(net195),
    .B(net385),
    .Y(_00199_));
 sky130_fd_sc_hd__xnor2_1 _06380_ (.A(_00198_),
    .B(_00199_),
    .Y(_00200_));
 sky130_fd_sc_hd__nand2b_1 _06381_ (.A_N(_00195_),
    .B(_00200_),
    .Y(_00201_));
 sky130_fd_sc_hd__xnor2_1 _06382_ (.A(_00195_),
    .B(_00200_),
    .Y(_00202_));
 sky130_fd_sc_hd__nand2b_1 _06383_ (.A_N(_00194_),
    .B(_00202_),
    .Y(_00203_));
 sky130_fd_sc_hd__xnor2_1 _06384_ (.A(_00194_),
    .B(_00202_),
    .Y(_00204_));
 sky130_fd_sc_hd__nand2_1 _06385_ (.A(net217),
    .B(net179),
    .Y(_00205_));
 sky130_fd_sc_hd__and4_1 _06386_ (.A(net241),
    .B(net232),
    .C(net171),
    .D(net163),
    .X(_00206_));
 sky130_fd_sc_hd__a22oi_1 _06387_ (.A1(net232),
    .A2(net171),
    .B1(net163),
    .B2(net241),
    .Y(_00207_));
 sky130_fd_sc_hd__nor2_1 _06388_ (.A(_00206_),
    .B(_00207_),
    .Y(_00208_));
 sky130_fd_sc_hd__xnor2_1 _06389_ (.A(_00205_),
    .B(_00208_),
    .Y(_00209_));
 sky130_fd_sc_hd__nand2_1 _06390_ (.A(net256),
    .B(net622),
    .Y(_00210_));
 sky130_fd_sc_hd__and4_1 _06391_ (.A(net438),
    .B(net346),
    .C(net614),
    .D(net597),
    .X(_00211_));
 sky130_fd_sc_hd__a22oi_2 _06392_ (.A1(net346),
    .A2(net614),
    .B1(net597),
    .B2(net438),
    .Y(_00212_));
 sky130_fd_sc_hd__or3_1 _06393_ (.A(_00210_),
    .B(_00211_),
    .C(_00212_),
    .X(_00213_));
 sky130_fd_sc_hd__o21ai_1 _06394_ (.A1(_00211_),
    .A2(_00212_),
    .B1(_00210_),
    .Y(_00214_));
 sky130_fd_sc_hd__o21bai_1 _06395_ (.A1(_00107_),
    .A2(_00109_),
    .B1_N(_00108_),
    .Y(_00215_));
 sky130_fd_sc_hd__nand3_1 _06396_ (.A(_00213_),
    .B(_00214_),
    .C(_00215_),
    .Y(_00216_));
 sky130_fd_sc_hd__a21o_1 _06397_ (.A1(_00213_),
    .A2(_00214_),
    .B1(_00215_),
    .X(_00217_));
 sky130_fd_sc_hd__nand3_1 _06398_ (.A(_00209_),
    .B(_00216_),
    .C(_00217_),
    .Y(_00218_));
 sky130_fd_sc_hd__a21o_1 _06399_ (.A1(_00216_),
    .A2(_00217_),
    .B1(_00209_),
    .X(_00219_));
 sky130_fd_sc_hd__a21bo_1 _06400_ (.A1(_00106_),
    .A2(_00114_),
    .B1_N(_00113_),
    .X(_00220_));
 sky130_fd_sc_hd__nand3_4 _06401_ (.A(_00218_),
    .B(_00219_),
    .C(_00220_),
    .Y(_00221_));
 sky130_fd_sc_hd__a21o_1 _06402_ (.A1(_00218_),
    .A2(_00219_),
    .B1(_00220_),
    .X(_00222_));
 sky130_fd_sc_hd__and3_1 _06403_ (.A(_00204_),
    .B(_00221_),
    .C(_00222_),
    .X(_00223_));
 sky130_fd_sc_hd__nand3_2 _06404_ (.A(_00204_),
    .B(_00221_),
    .C(_00222_),
    .Y(_00224_));
 sky130_fd_sc_hd__a21oi_2 _06405_ (.A1(_00221_),
    .A2(_00222_),
    .B1(_00204_),
    .Y(_00225_));
 sky130_fd_sc_hd__a211oi_4 _06406_ (.A1(_00118_),
    .A2(_00121_),
    .B1(_00223_),
    .C1(_00225_),
    .Y(_00226_));
 sky130_fd_sc_hd__o211a_1 _06407_ (.A1(_00223_),
    .A2(_00225_),
    .B1(_00118_),
    .C1(_00121_),
    .X(_00227_));
 sky130_fd_sc_hd__nor4_1 _06408_ (.A(_00191_),
    .B(_00193_),
    .C(_00226_),
    .D(_00227_),
    .Y(_00228_));
 sky130_fd_sc_hd__or4_2 _06409_ (.A(_00191_),
    .B(_00193_),
    .C(_00226_),
    .D(_00227_),
    .X(_00229_));
 sky130_fd_sc_hd__o22ai_2 _06410_ (.A1(_00191_),
    .A2(_00193_),
    .B1(_00226_),
    .B2(_00227_),
    .Y(_00230_));
 sky130_fd_sc_hd__o211ai_4 _06411_ (.A1(_00123_),
    .A2(net150),
    .B1(_00229_),
    .C1(_00230_),
    .Y(_00231_));
 sky130_fd_sc_hd__a211o_1 _06412_ (.A1(_00229_),
    .A2(_00230_),
    .B1(_00123_),
    .C1(_00125_),
    .X(_00232_));
 sky130_fd_sc_hd__and4bb_1 _06413_ (.A_N(_00172_),
    .B_N(_00173_),
    .C(_00231_),
    .D(_00232_),
    .X(_00233_));
 sky130_fd_sc_hd__or4bb_1 _06414_ (.A(_00172_),
    .B(_00173_),
    .C_N(_00231_),
    .D_N(_00232_),
    .X(_00234_));
 sky130_fd_sc_hd__a2bb2oi_1 _06415_ (.A1_N(_00172_),
    .A2_N(_00173_),
    .B1(_00231_),
    .B2(_00232_),
    .Y(_00235_));
 sky130_fd_sc_hd__a211oi_2 _06416_ (.A1(_00128_),
    .A2(_00130_),
    .B1(_00233_),
    .C1(_00235_),
    .Y(_00236_));
 sky130_fd_sc_hd__o211a_1 _06417_ (.A1(_00233_),
    .A2(_00235_),
    .B1(_00128_),
    .C1(_00130_),
    .X(_00237_));
 sky130_fd_sc_hd__nor2_1 _06418_ (.A(_00236_),
    .B(_00237_),
    .Y(_00238_));
 sky130_fd_sc_hd__and2b_1 _06419_ (.A_N(_00144_),
    .B(_00238_),
    .X(_00239_));
 sky130_fd_sc_hd__xnor2_1 _06420_ (.A(_00144_),
    .B(_00238_),
    .Y(_00240_));
 sky130_fd_sc_hd__a32oi_2 _06421_ (.A1(_00130_),
    .A2(_00131_),
    .A3(_00133_),
    .B1(_00134_),
    .B2(_00045_),
    .Y(_00241_));
 sky130_fd_sc_hd__and2b_1 _06422_ (.A_N(_00241_),
    .B(_00240_),
    .X(_00242_));
 sky130_fd_sc_hd__inv_2 _06423_ (.A(_00242_),
    .Y(_00243_));
 sky130_fd_sc_hd__xnor2_1 _06424_ (.A(_00240_),
    .B(_00241_),
    .Y(_00244_));
 sky130_fd_sc_hd__and2b_1 _06425_ (.A_N(_00137_),
    .B(_00244_),
    .X(_00245_));
 sky130_fd_sc_hd__xnor2_1 _06426_ (.A(_00137_),
    .B(_00244_),
    .Y(_00246_));
 sky130_fd_sc_hd__and2_1 _06427_ (.A(_00139_),
    .B(_00246_),
    .X(_00247_));
 sky130_fd_sc_hd__xor2_1 _06428_ (.A(_00139_),
    .B(_00246_),
    .X(_00248_));
 sky130_fd_sc_hd__inv_2 _06429_ (.A(_00248_),
    .Y(_00249_));
 sky130_fd_sc_hd__and2_1 _06430_ (.A(_00038_),
    .B(_00142_),
    .X(_00250_));
 sky130_fd_sc_hd__o21a_1 _06431_ (.A1(_00034_),
    .A2(_00036_),
    .B1(_00141_),
    .X(_00251_));
 sky130_fd_sc_hd__a31o_1 _06432_ (.A1(_00038_),
    .A2(_00040_),
    .A3(_00142_),
    .B1(_00251_),
    .X(_00252_));
 sky130_fd_sc_hd__and3b_1 _06433_ (.A_N(_05070_),
    .B(_00041_),
    .C(_00250_),
    .X(_00253_));
 sky130_fd_sc_hd__nor2_1 _06434_ (.A(_00252_),
    .B(_00253_),
    .Y(_00254_));
 sky130_fd_sc_hd__nor2_1 _06435_ (.A(_00249_),
    .B(_00254_),
    .Y(_00255_));
 sky130_fd_sc_hd__xnor2_1 _06436_ (.A(_00248_),
    .B(_00254_),
    .Y(net77));
 sky130_fd_sc_hd__o21ai_1 _06437_ (.A1(_00170_),
    .A2(_00172_),
    .B1(_00150_),
    .Y(_00256_));
 sky130_fd_sc_hd__or3_1 _06438_ (.A(_00150_),
    .B(_00170_),
    .C(_00172_),
    .X(_00257_));
 sky130_fd_sc_hd__and2_1 _06439_ (.A(_00256_),
    .B(_00257_),
    .X(_00258_));
 sky130_fd_sc_hd__and4_1 _06440_ (.A(net498),
    .B(net518),
    .C(net363),
    .D(net355),
    .X(_00259_));
 sky130_fd_sc_hd__a22o_1 _06441_ (.A1(net498),
    .A2(net363),
    .B1(net355),
    .B2(net518),
    .X(_00260_));
 sky130_fd_sc_hd__and2b_1 _06442_ (.A_N(_00259_),
    .B(_00260_),
    .X(_00261_));
 sky130_fd_sc_hd__nand2_1 _06443_ (.A(net604),
    .B(net338),
    .Y(_00262_));
 sky130_fd_sc_hd__xnor2_1 _06444_ (.A(_00261_),
    .B(_00262_),
    .Y(_00263_));
 sky130_fd_sc_hd__a31oi_2 _06445_ (.A1(net629),
    .A2(net338),
    .A3(_00147_),
    .B1(_00145_),
    .Y(_00264_));
 sky130_fd_sc_hd__and2b_1 _06446_ (.A_N(_00264_),
    .B(_00263_),
    .X(_00265_));
 sky130_fd_sc_hd__xnor2_1 _06447_ (.A(_00263_),
    .B(_00264_),
    .Y(_00266_));
 sky130_fd_sc_hd__nand2_1 _06448_ (.A(net629),
    .B(net333),
    .Y(_00267_));
 sky130_fd_sc_hd__xor2_1 _06449_ (.A(_00266_),
    .B(_00267_),
    .X(_00268_));
 sky130_fd_sc_hd__a31o_1 _06450_ (.A1(net499),
    .A2(net371),
    .A3(_00157_),
    .B1(_00155_),
    .X(_00269_));
 sky130_fd_sc_hd__o21ba_1 _06451_ (.A1(_00174_),
    .A2(_00176_),
    .B1_N(_00175_),
    .X(_00270_));
 sky130_fd_sc_hd__and4_1 _06452_ (.A(net483),
    .B(net475),
    .C(net395),
    .D(net379),
    .X(_00271_));
 sky130_fd_sc_hd__a22oi_1 _06453_ (.A1(net475),
    .A2(net395),
    .B1(net379),
    .B2(net483),
    .Y(_00272_));
 sky130_fd_sc_hd__nor2_1 _06454_ (.A(_00271_),
    .B(_00272_),
    .Y(_00273_));
 sky130_fd_sc_hd__nand2_1 _06455_ (.A(net491),
    .B(net371),
    .Y(_00274_));
 sky130_fd_sc_hd__xnor2_1 _06456_ (.A(_00273_),
    .B(_00274_),
    .Y(_00275_));
 sky130_fd_sc_hd__nand2b_1 _06457_ (.A_N(_00270_),
    .B(_00275_),
    .Y(_00276_));
 sky130_fd_sc_hd__xnor2_1 _06458_ (.A(_00270_),
    .B(_00275_),
    .Y(_00277_));
 sky130_fd_sc_hd__nand2_1 _06459_ (.A(_00269_),
    .B(_00277_),
    .Y(_00278_));
 sky130_fd_sc_hd__xnor2_1 _06460_ (.A(_00269_),
    .B(_00277_),
    .Y(_00279_));
 sky130_fd_sc_hd__a21oi_2 _06461_ (.A1(_00160_),
    .A2(_00162_),
    .B1(_00279_),
    .Y(_00280_));
 sky130_fd_sc_hd__inv_2 _06462_ (.A(_00280_),
    .Y(_00281_));
 sky130_fd_sc_hd__and3_1 _06463_ (.A(_00160_),
    .B(_00162_),
    .C(_00279_),
    .X(_00282_));
 sky130_fd_sc_hd__nor3_1 _06464_ (.A(_00268_),
    .B(_00280_),
    .C(_00282_),
    .Y(_00283_));
 sky130_fd_sc_hd__or3_1 _06465_ (.A(_00268_),
    .B(_00280_),
    .C(_00282_),
    .X(_00284_));
 sky130_fd_sc_hd__o21a_1 _06466_ (.A1(_00280_),
    .A2(_00282_),
    .B1(_00268_),
    .X(_00285_));
 sky130_fd_sc_hd__a211oi_2 _06467_ (.A1(_00189_),
    .A2(_00192_),
    .B1(_00283_),
    .C1(_00285_),
    .Y(_00286_));
 sky130_fd_sc_hd__o211a_1 _06468_ (.A1(_00283_),
    .A2(_00285_),
    .B1(_00189_),
    .C1(_00192_),
    .X(_00288_));
 sky130_fd_sc_hd__a211oi_2 _06469_ (.A1(_00165_),
    .A2(_00168_),
    .B1(_00286_),
    .C1(_00288_),
    .Y(_00289_));
 sky130_fd_sc_hd__o211a_1 _06470_ (.A1(_00286_),
    .A2(_00288_),
    .B1(_00165_),
    .C1(_00168_),
    .X(_00290_));
 sky130_fd_sc_hd__and4_1 _06471_ (.A(net453),
    .B(net447),
    .C(net418),
    .D(net410),
    .X(_00291_));
 sky130_fd_sc_hd__a22oi_1 _06472_ (.A1(net448),
    .A2(net418),
    .B1(net410),
    .B2(net454),
    .Y(_00292_));
 sky130_fd_sc_hd__nor2_1 _06473_ (.A(_00291_),
    .B(_00292_),
    .Y(_00293_));
 sky130_fd_sc_hd__nand2_1 _06474_ (.A(net460),
    .B(net402),
    .Y(_00294_));
 sky130_fd_sc_hd__xnor2_1 _06475_ (.A(_00293_),
    .B(_00294_),
    .Y(_00295_));
 sky130_fd_sc_hd__and4_1 _06476_ (.A(net189),
    .B(net432),
    .C(net467),
    .D(net386),
    .X(_00296_));
 sky130_fd_sc_hd__a22oi_1 _06477_ (.A1(net432),
    .A2(net467),
    .B1(net386),
    .B2(net189),
    .Y(_00297_));
 sky130_fd_sc_hd__nor2_1 _06478_ (.A(_00296_),
    .B(_00297_),
    .Y(_00299_));
 sky130_fd_sc_hd__nand2_1 _06479_ (.A(net549),
    .B(net424),
    .Y(_00300_));
 sky130_fd_sc_hd__xnor2_1 _06480_ (.A(_00299_),
    .B(_00300_),
    .Y(_00301_));
 sky130_fd_sc_hd__o21ba_1 _06481_ (.A1(_00179_),
    .A2(_00181_),
    .B1_N(_00180_),
    .X(_00302_));
 sky130_fd_sc_hd__and2b_1 _06482_ (.A_N(_00302_),
    .B(_00301_),
    .X(_00303_));
 sky130_fd_sc_hd__xnor2_1 _06483_ (.A(_00301_),
    .B(_00302_),
    .Y(_00304_));
 sky130_fd_sc_hd__and2_1 _06484_ (.A(_00295_),
    .B(_00304_),
    .X(_00305_));
 sky130_fd_sc_hd__xnor2_1 _06485_ (.A(_00295_),
    .B(_00304_),
    .Y(_00306_));
 sky130_fd_sc_hd__a21o_1 _06486_ (.A1(_00201_),
    .A2(_00203_),
    .B1(_00306_),
    .X(_00307_));
 sky130_fd_sc_hd__inv_2 _06487_ (.A(_00307_),
    .Y(_00308_));
 sky130_fd_sc_hd__nand3_1 _06488_ (.A(_00201_),
    .B(_00203_),
    .C(_00306_),
    .Y(_00310_));
 sky130_fd_sc_hd__o211a_1 _06489_ (.A1(_00185_),
    .A2(_00187_),
    .B1(_00307_),
    .C1(_00310_),
    .X(_00311_));
 sky130_fd_sc_hd__a211oi_2 _06490_ (.A1(_00307_),
    .A2(_00310_),
    .B1(_00185_),
    .C1(_00187_),
    .Y(_00312_));
 sky130_fd_sc_hd__o21ba_1 _06491_ (.A1(_00197_),
    .A2(_00199_),
    .B1_N(_00196_),
    .X(_00313_));
 sky130_fd_sc_hd__o21ba_1 _06492_ (.A1(_00205_),
    .A2(_00207_),
    .B1_N(_00206_),
    .X(_00314_));
 sky130_fd_sc_hd__and4_1 _06493_ (.A(net213),
    .B(net204),
    .C(net224),
    .D(net179),
    .X(_00315_));
 sky130_fd_sc_hd__a22oi_1 _06494_ (.A1(net204),
    .A2(net224),
    .B1(net179),
    .B2(net213),
    .Y(_00316_));
 sky130_fd_sc_hd__nor2_1 _06495_ (.A(_00315_),
    .B(_00316_),
    .Y(_00317_));
 sky130_fd_sc_hd__nand2_1 _06496_ (.A(net195),
    .B(net300),
    .Y(_00318_));
 sky130_fd_sc_hd__xnor2_1 _06497_ (.A(_00317_),
    .B(_00318_),
    .Y(_00319_));
 sky130_fd_sc_hd__nand2b_1 _06498_ (.A_N(_00314_),
    .B(_00319_),
    .Y(_00321_));
 sky130_fd_sc_hd__xnor2_1 _06499_ (.A(_00314_),
    .B(_00319_),
    .Y(_00322_));
 sky130_fd_sc_hd__nand2b_1 _06500_ (.A_N(_00313_),
    .B(_00322_),
    .Y(_00323_));
 sky130_fd_sc_hd__xnor2_1 _06501_ (.A(_00313_),
    .B(_00322_),
    .Y(_00324_));
 sky130_fd_sc_hd__nand2_1 _06502_ (.A(net217),
    .B(net171),
    .Y(_00325_));
 sky130_fd_sc_hd__and4_1 _06503_ (.A(net241),
    .B(net232),
    .C(net163),
    .D(net620),
    .X(_00326_));
 sky130_fd_sc_hd__a22oi_1 _06504_ (.A1(net234),
    .A2(net163),
    .B1(net620),
    .B2(net241),
    .Y(_00327_));
 sky130_fd_sc_hd__nor2_1 _06505_ (.A(_00326_),
    .B(_00327_),
    .Y(_00328_));
 sky130_fd_sc_hd__xnor2_1 _06506_ (.A(_00325_),
    .B(_00328_),
    .Y(_00329_));
 sky130_fd_sc_hd__nand2_1 _06507_ (.A(net256),
    .B(net614),
    .Y(_00330_));
 sky130_fd_sc_hd__and4_1 _06508_ (.A(net438),
    .B(net346),
    .C(net597),
    .D(net589),
    .X(_00332_));
 sky130_fd_sc_hd__a22oi_2 _06509_ (.A1(net346),
    .A2(net597),
    .B1(net589),
    .B2(net438),
    .Y(_00333_));
 sky130_fd_sc_hd__or3_1 _06510_ (.A(_00330_),
    .B(_00332_),
    .C(_00333_),
    .X(_00334_));
 sky130_fd_sc_hd__o21ai_1 _06511_ (.A1(_00332_),
    .A2(_00333_),
    .B1(_00330_),
    .Y(_00335_));
 sky130_fd_sc_hd__o21bai_1 _06512_ (.A1(_00210_),
    .A2(_00212_),
    .B1_N(_00211_),
    .Y(_00336_));
 sky130_fd_sc_hd__nand3_1 _06513_ (.A(_00334_),
    .B(_00335_),
    .C(_00336_),
    .Y(_00337_));
 sky130_fd_sc_hd__a21o_1 _06514_ (.A1(_00334_),
    .A2(_00335_),
    .B1(_00336_),
    .X(_00338_));
 sky130_fd_sc_hd__nand3_1 _06515_ (.A(_00329_),
    .B(_00337_),
    .C(_00338_),
    .Y(_00339_));
 sky130_fd_sc_hd__a21o_1 _06516_ (.A1(_00337_),
    .A2(_00338_),
    .B1(_00329_),
    .X(_00340_));
 sky130_fd_sc_hd__a21bo_1 _06517_ (.A1(_00209_),
    .A2(_00217_),
    .B1_N(_00216_),
    .X(_00341_));
 sky130_fd_sc_hd__nand3_4 _06518_ (.A(_00339_),
    .B(_00340_),
    .C(_00341_),
    .Y(_00343_));
 sky130_fd_sc_hd__a21o_1 _06519_ (.A1(_00339_),
    .A2(_00340_),
    .B1(_00341_),
    .X(_00344_));
 sky130_fd_sc_hd__and3_1 _06520_ (.A(_00324_),
    .B(_00343_),
    .C(_00344_),
    .X(_00345_));
 sky130_fd_sc_hd__nand3_2 _06521_ (.A(_00324_),
    .B(_00343_),
    .C(_00344_),
    .Y(_00346_));
 sky130_fd_sc_hd__a21oi_2 _06522_ (.A1(_00343_),
    .A2(_00344_),
    .B1(_00324_),
    .Y(_00347_));
 sky130_fd_sc_hd__a211oi_4 _06523_ (.A1(_00221_),
    .A2(_00224_),
    .B1(_00345_),
    .C1(_00347_),
    .Y(_00348_));
 sky130_fd_sc_hd__o211a_1 _06524_ (.A1(_00345_),
    .A2(_00347_),
    .B1(_00221_),
    .C1(_00224_),
    .X(_00349_));
 sky130_fd_sc_hd__nor4_1 _06525_ (.A(_00311_),
    .B(_00312_),
    .C(_00348_),
    .D(_00349_),
    .Y(_00350_));
 sky130_fd_sc_hd__or4_2 _06526_ (.A(_00311_),
    .B(_00312_),
    .C(_00348_),
    .D(_00349_),
    .X(_00351_));
 sky130_fd_sc_hd__o22ai_2 _06527_ (.A1(_00311_),
    .A2(_00312_),
    .B1(_00348_),
    .B2(_00349_),
    .Y(_00352_));
 sky130_fd_sc_hd__o211ai_4 _06528_ (.A1(_00226_),
    .A2(net149),
    .B1(_00351_),
    .C1(_00352_),
    .Y(_00354_));
 sky130_fd_sc_hd__a211o_1 _06529_ (.A1(_00351_),
    .A2(_00352_),
    .B1(_00226_),
    .C1(_00228_),
    .X(_00355_));
 sky130_fd_sc_hd__and4bb_1 _06530_ (.A_N(_00289_),
    .B_N(_00290_),
    .C(_00354_),
    .D(_00355_),
    .X(_00356_));
 sky130_fd_sc_hd__or4bb_1 _06531_ (.A(_00289_),
    .B(_00290_),
    .C_N(_00354_),
    .D_N(_00355_),
    .X(_00357_));
 sky130_fd_sc_hd__a2bb2oi_1 _06532_ (.A1_N(_00289_),
    .A2_N(_00290_),
    .B1(_00354_),
    .B2(_00355_),
    .Y(_00358_));
 sky130_fd_sc_hd__a211o_1 _06533_ (.A1(_00231_),
    .A2(_00234_),
    .B1(_00356_),
    .C1(_00358_),
    .X(_00359_));
 sky130_fd_sc_hd__o211ai_2 _06534_ (.A1(_00356_),
    .A2(_00358_),
    .B1(_00231_),
    .C1(_00234_),
    .Y(_00360_));
 sky130_fd_sc_hd__nand3_2 _06535_ (.A(_00258_),
    .B(_00359_),
    .C(_00360_),
    .Y(_00361_));
 sky130_fd_sc_hd__a21o_1 _06536_ (.A1(_00359_),
    .A2(_00360_),
    .B1(_00258_),
    .X(_00362_));
 sky130_fd_sc_hd__o211ai_2 _06537_ (.A1(_00236_),
    .A2(_00239_),
    .B1(_00361_),
    .C1(_00362_),
    .Y(_00363_));
 sky130_fd_sc_hd__a211o_1 _06538_ (.A1(_00361_),
    .A2(_00362_),
    .B1(_00236_),
    .C1(_00239_),
    .X(_00365_));
 sky130_fd_sc_hd__nand2_1 _06539_ (.A(_00363_),
    .B(_00365_),
    .Y(_00366_));
 sky130_fd_sc_hd__nor2_1 _06540_ (.A(_00243_),
    .B(_00366_),
    .Y(_00367_));
 sky130_fd_sc_hd__xnor2_1 _06541_ (.A(_00242_),
    .B(_00366_),
    .Y(_00368_));
 sky130_fd_sc_hd__xor2_1 _06542_ (.A(_00245_),
    .B(_00368_),
    .X(_00369_));
 sky130_fd_sc_hd__nor2_1 _06543_ (.A(_00247_),
    .B(_00255_),
    .Y(_00370_));
 sky130_fd_sc_hd__xnor2_1 _06544_ (.A(_00369_),
    .B(_00370_),
    .Y(net78));
 sky130_fd_sc_hd__a31oi_1 _06545_ (.A1(net629),
    .A2(net333),
    .A3(_00266_),
    .B1(_00265_),
    .Y(_00371_));
 sky130_fd_sc_hd__o21ba_1 _06546_ (.A1(_00286_),
    .A2(_00289_),
    .B1_N(_00371_),
    .X(_00372_));
 sky130_fd_sc_hd__or3b_1 _06547_ (.A(_00286_),
    .B(_00289_),
    .C_N(_00371_),
    .X(_00373_));
 sky130_fd_sc_hd__and2b_1 _06548_ (.A_N(_00372_),
    .B(_00373_),
    .X(_00375_));
 sky130_fd_sc_hd__a22o_1 _06549_ (.A1(net604),
    .A2(net332),
    .B1(net325),
    .B2(net629),
    .X(_00376_));
 sky130_fd_sc_hd__nand4_2 _06550_ (.A(net604),
    .B(net630),
    .C(net332),
    .D(net325),
    .Y(_00377_));
 sky130_fd_sc_hd__and4_1 _06551_ (.A(net490),
    .B(net498),
    .C(net363),
    .D(net355),
    .X(_00378_));
 sky130_fd_sc_hd__a22o_1 _06552_ (.A1(net490),
    .A2(net363),
    .B1(net355),
    .B2(net498),
    .X(_00379_));
 sky130_fd_sc_hd__and2b_1 _06553_ (.A_N(_00378_),
    .B(_00379_),
    .X(_00380_));
 sky130_fd_sc_hd__nand2_1 _06554_ (.A(net518),
    .B(net338),
    .Y(_00381_));
 sky130_fd_sc_hd__xnor2_1 _06555_ (.A(_00380_),
    .B(_00381_),
    .Y(_00382_));
 sky130_fd_sc_hd__a31o_1 _06556_ (.A1(net604),
    .A2(net338),
    .A3(_00260_),
    .B1(_00259_),
    .X(_00383_));
 sky130_fd_sc_hd__nand2_1 _06557_ (.A(_00382_),
    .B(_00383_),
    .Y(_00384_));
 sky130_fd_sc_hd__or2_1 _06558_ (.A(_00382_),
    .B(_00383_),
    .X(_00386_));
 sky130_fd_sc_hd__nand4_2 _06559_ (.A(_00376_),
    .B(_00377_),
    .C(_00384_),
    .D(_00386_),
    .Y(_00387_));
 sky130_fd_sc_hd__a22o_1 _06560_ (.A1(_00376_),
    .A2(_00377_),
    .B1(_00384_),
    .B2(_00386_),
    .X(_00388_));
 sky130_fd_sc_hd__a31o_1 _06561_ (.A1(net491),
    .A2(net371),
    .A3(_00273_),
    .B1(_00271_),
    .X(_00389_));
 sky130_fd_sc_hd__o21ba_1 _06562_ (.A1(_00292_),
    .A2(_00294_),
    .B1_N(_00291_),
    .X(_00390_));
 sky130_fd_sc_hd__and4_1 _06563_ (.A(net475),
    .B(net460),
    .C(net395),
    .D(net379),
    .X(_00391_));
 sky130_fd_sc_hd__a22oi_1 _06564_ (.A1(net460),
    .A2(net395),
    .B1(net379),
    .B2(net475),
    .Y(_00392_));
 sky130_fd_sc_hd__nor2_1 _06565_ (.A(_00391_),
    .B(_00392_),
    .Y(_00393_));
 sky130_fd_sc_hd__nand2_1 _06566_ (.A(net483),
    .B(net371),
    .Y(_00394_));
 sky130_fd_sc_hd__xnor2_1 _06567_ (.A(_00393_),
    .B(_00394_),
    .Y(_00395_));
 sky130_fd_sc_hd__nand2b_1 _06568_ (.A_N(_00390_),
    .B(_00395_),
    .Y(_00397_));
 sky130_fd_sc_hd__xnor2_1 _06569_ (.A(_00390_),
    .B(_00395_),
    .Y(_00398_));
 sky130_fd_sc_hd__nand2_1 _06570_ (.A(_00389_),
    .B(_00398_),
    .Y(_00399_));
 sky130_fd_sc_hd__xnor2_1 _06571_ (.A(_00389_),
    .B(_00398_),
    .Y(_00400_));
 sky130_fd_sc_hd__a21o_1 _06572_ (.A1(_00276_),
    .A2(_00278_),
    .B1(_00400_),
    .X(_00401_));
 sky130_fd_sc_hd__nand3_1 _06573_ (.A(_00276_),
    .B(_00278_),
    .C(_00400_),
    .Y(_00402_));
 sky130_fd_sc_hd__nand4_2 _06574_ (.A(_00387_),
    .B(_00388_),
    .C(_00401_),
    .D(_00402_),
    .Y(_00403_));
 sky130_fd_sc_hd__a22o_1 _06575_ (.A1(_00387_),
    .A2(_00388_),
    .B1(_00401_),
    .B2(_00402_),
    .X(_00404_));
 sky130_fd_sc_hd__o211a_1 _06576_ (.A1(_00308_),
    .A2(_00311_),
    .B1(_00403_),
    .C1(_00404_),
    .X(_00405_));
 sky130_fd_sc_hd__a211oi_1 _06577_ (.A1(_00403_),
    .A2(_00404_),
    .B1(_00308_),
    .C1(_00311_),
    .Y(_00406_));
 sky130_fd_sc_hd__a211oi_1 _06578_ (.A1(_00281_),
    .A2(_00284_),
    .B1(_00405_),
    .C1(_00406_),
    .Y(_00408_));
 sky130_fd_sc_hd__o211a_1 _06579_ (.A1(_00405_),
    .A2(_00406_),
    .B1(_00281_),
    .C1(_00284_),
    .X(_00409_));
 sky130_fd_sc_hd__and4_1 _06580_ (.A(net549),
    .B(net448),
    .C(net417),
    .D(net409),
    .X(_00410_));
 sky130_fd_sc_hd__a22oi_1 _06581_ (.A1(net549),
    .A2(net417),
    .B1(net409),
    .B2(net448),
    .Y(_00411_));
 sky130_fd_sc_hd__nor2_1 _06582_ (.A(_00410_),
    .B(_00411_),
    .Y(_00412_));
 sky130_fd_sc_hd__nand2_1 _06583_ (.A(net454),
    .B(net403),
    .Y(_00413_));
 sky130_fd_sc_hd__xnor2_1 _06584_ (.A(_00412_),
    .B(_00413_),
    .Y(_00414_));
 sky130_fd_sc_hd__and4_1 _06585_ (.A(net189),
    .B(net432),
    .C(net386),
    .D(net300),
    .X(_00415_));
 sky130_fd_sc_hd__a22o_1 _06586_ (.A1(net432),
    .A2(net387),
    .B1(net300),
    .B2(net189),
    .X(_00416_));
 sky130_fd_sc_hd__and2b_1 _06587_ (.A_N(_00415_),
    .B(_00416_),
    .X(_00417_));
 sky130_fd_sc_hd__nand2_1 _06588_ (.A(net467),
    .B(net424),
    .Y(_00419_));
 sky130_fd_sc_hd__xnor2_1 _06589_ (.A(_00417_),
    .B(_00419_),
    .Y(_00420_));
 sky130_fd_sc_hd__o21ba_1 _06590_ (.A1(_00297_),
    .A2(_00300_),
    .B1_N(_00296_),
    .X(_00421_));
 sky130_fd_sc_hd__and2b_1 _06591_ (.A_N(_00421_),
    .B(_00420_),
    .X(_00422_));
 sky130_fd_sc_hd__xnor2_1 _06592_ (.A(_00420_),
    .B(_00421_),
    .Y(_00423_));
 sky130_fd_sc_hd__and2_1 _06593_ (.A(_00414_),
    .B(_00423_),
    .X(_00424_));
 sky130_fd_sc_hd__xnor2_1 _06594_ (.A(_00414_),
    .B(_00423_),
    .Y(_00425_));
 sky130_fd_sc_hd__a21o_1 _06595_ (.A1(_00321_),
    .A2(_00323_),
    .B1(_00425_),
    .X(_00426_));
 sky130_fd_sc_hd__nand3_2 _06596_ (.A(_00321_),
    .B(_00323_),
    .C(_00425_),
    .Y(_00427_));
 sky130_fd_sc_hd__o211a_1 _06597_ (.A1(_00303_),
    .A2(_00305_),
    .B1(_00426_),
    .C1(_00427_),
    .X(_00428_));
 sky130_fd_sc_hd__o211ai_2 _06598_ (.A1(_00303_),
    .A2(_00305_),
    .B1(_00426_),
    .C1(_00427_),
    .Y(_00430_));
 sky130_fd_sc_hd__a211oi_2 _06599_ (.A1(_00426_),
    .A2(_00427_),
    .B1(_00303_),
    .C1(_00305_),
    .Y(_00431_));
 sky130_fd_sc_hd__a31o_1 _06600_ (.A1(net197),
    .A2(net300),
    .A3(_00317_),
    .B1(_00315_),
    .X(_00432_));
 sky130_fd_sc_hd__o21bai_1 _06601_ (.A1(_00325_),
    .A2(_00327_),
    .B1_N(_00326_),
    .Y(_00433_));
 sky130_fd_sc_hd__nand4_1 _06602_ (.A(net213),
    .B(net204),
    .C(net179),
    .D(net171),
    .Y(_00434_));
 sky130_fd_sc_hd__a22o_1 _06603_ (.A1(net204),
    .A2(net179),
    .B1(net171),
    .B2(net213),
    .X(_00435_));
 sky130_fd_sc_hd__nand2_1 _06604_ (.A(net197),
    .B(net224),
    .Y(_00436_));
 sky130_fd_sc_hd__nand3b_1 _06605_ (.A_N(_00436_),
    .B(_00435_),
    .C(_00434_),
    .Y(_00437_));
 sky130_fd_sc_hd__a21bo_1 _06606_ (.A1(_00434_),
    .A2(_00435_),
    .B1_N(_00436_),
    .X(_00438_));
 sky130_fd_sc_hd__and3_1 _06607_ (.A(_00433_),
    .B(_00437_),
    .C(_00438_),
    .X(_00439_));
 sky130_fd_sc_hd__a21o_1 _06608_ (.A1(_00437_),
    .A2(_00438_),
    .B1(_00433_),
    .X(_00441_));
 sky130_fd_sc_hd__and2b_1 _06609_ (.A_N(_00439_),
    .B(_00441_),
    .X(_00442_));
 sky130_fd_sc_hd__xor2_2 _06610_ (.A(_00432_),
    .B(_00442_),
    .X(_00443_));
 sky130_fd_sc_hd__nand2_1 _06611_ (.A(net217),
    .B(net163),
    .Y(_00444_));
 sky130_fd_sc_hd__and4_1 _06612_ (.A(net240),
    .B(net233),
    .C(net620),
    .D(net612),
    .X(_00445_));
 sky130_fd_sc_hd__a22oi_1 _06613_ (.A1(net233),
    .A2(net620),
    .B1(net612),
    .B2(net240),
    .Y(_00446_));
 sky130_fd_sc_hd__nor2_1 _06614_ (.A(_00445_),
    .B(_00446_),
    .Y(_00447_));
 sky130_fd_sc_hd__xnor2_1 _06615_ (.A(_00444_),
    .B(_00447_),
    .Y(_00448_));
 sky130_fd_sc_hd__nand2_1 _06616_ (.A(net258),
    .B(net597),
    .Y(_00449_));
 sky130_fd_sc_hd__and4_1 _06617_ (.A(net438),
    .B(net346),
    .C(net589),
    .D(net581),
    .X(_00450_));
 sky130_fd_sc_hd__a22oi_2 _06618_ (.A1(net348),
    .A2(net589),
    .B1(net581),
    .B2(net438),
    .Y(_00452_));
 sky130_fd_sc_hd__or3_1 _06619_ (.A(_00449_),
    .B(_00450_),
    .C(_00452_),
    .X(_00453_));
 sky130_fd_sc_hd__o21ai_1 _06620_ (.A1(_00450_),
    .A2(_00452_),
    .B1(_00449_),
    .Y(_00454_));
 sky130_fd_sc_hd__o21bai_1 _06621_ (.A1(_00330_),
    .A2(_00333_),
    .B1_N(_00332_),
    .Y(_00455_));
 sky130_fd_sc_hd__nand3_1 _06622_ (.A(_00453_),
    .B(_00454_),
    .C(_00455_),
    .Y(_00456_));
 sky130_fd_sc_hd__a21o_1 _06623_ (.A1(_00453_),
    .A2(_00454_),
    .B1(_00455_),
    .X(_00457_));
 sky130_fd_sc_hd__nand3_2 _06624_ (.A(_00448_),
    .B(_00456_),
    .C(_00457_),
    .Y(_00458_));
 sky130_fd_sc_hd__a21o_1 _06625_ (.A1(_00456_),
    .A2(_00457_),
    .B1(_00448_),
    .X(_00459_));
 sky130_fd_sc_hd__a21bo_1 _06626_ (.A1(_00329_),
    .A2(_00338_),
    .B1_N(_00337_),
    .X(_00460_));
 sky130_fd_sc_hd__nand3_4 _06627_ (.A(_00458_),
    .B(_00459_),
    .C(_00460_),
    .Y(_00461_));
 sky130_fd_sc_hd__a21o_1 _06628_ (.A1(_00458_),
    .A2(_00459_),
    .B1(_00460_),
    .X(_00463_));
 sky130_fd_sc_hd__and3_1 _06629_ (.A(_00443_),
    .B(_00461_),
    .C(_00463_),
    .X(_00464_));
 sky130_fd_sc_hd__nand3_2 _06630_ (.A(_00443_),
    .B(_00461_),
    .C(_00463_),
    .Y(_00465_));
 sky130_fd_sc_hd__a21oi_2 _06631_ (.A1(_00461_),
    .A2(_00463_),
    .B1(_00443_),
    .Y(_00466_));
 sky130_fd_sc_hd__a211oi_4 _06632_ (.A1(_00343_),
    .A2(_00346_),
    .B1(_00464_),
    .C1(_00466_),
    .Y(_00467_));
 sky130_fd_sc_hd__o211a_1 _06633_ (.A1(_00464_),
    .A2(_00466_),
    .B1(_00343_),
    .C1(_00346_),
    .X(_00468_));
 sky130_fd_sc_hd__nor4_1 _06634_ (.A(_00428_),
    .B(_00431_),
    .C(_00467_),
    .D(_00468_),
    .Y(_00469_));
 sky130_fd_sc_hd__or4_2 _06635_ (.A(_00428_),
    .B(_00431_),
    .C(_00467_),
    .D(_00468_),
    .X(_00470_));
 sky130_fd_sc_hd__o22ai_2 _06636_ (.A1(_00428_),
    .A2(_00431_),
    .B1(_00467_),
    .B2(_00468_),
    .Y(_00471_));
 sky130_fd_sc_hd__o211ai_4 _06637_ (.A1(_00348_),
    .A2(net148),
    .B1(_00470_),
    .C1(_00471_),
    .Y(_00472_));
 sky130_fd_sc_hd__a211o_1 _06638_ (.A1(_00470_),
    .A2(_00471_),
    .B1(_00348_),
    .C1(_00350_),
    .X(_00474_));
 sky130_fd_sc_hd__and4bb_1 _06639_ (.A_N(_00408_),
    .B_N(_00409_),
    .C(_00472_),
    .D(_00474_),
    .X(_00475_));
 sky130_fd_sc_hd__or4bb_1 _06640_ (.A(_00408_),
    .B(_00409_),
    .C_N(_00472_),
    .D_N(_00474_),
    .X(_00476_));
 sky130_fd_sc_hd__a2bb2oi_1 _06641_ (.A1_N(_00408_),
    .A2_N(_00409_),
    .B1(_00472_),
    .B2(_00474_),
    .Y(_00477_));
 sky130_fd_sc_hd__a211o_1 _06642_ (.A1(_00354_),
    .A2(_00357_),
    .B1(_00475_),
    .C1(_00477_),
    .X(_00478_));
 sky130_fd_sc_hd__o211ai_1 _06643_ (.A1(_00475_),
    .A2(_00477_),
    .B1(_00354_),
    .C1(_00357_),
    .Y(_00479_));
 sky130_fd_sc_hd__and3_1 _06644_ (.A(_00375_),
    .B(_00478_),
    .C(_00479_),
    .X(_00480_));
 sky130_fd_sc_hd__nand3_1 _06645_ (.A(_00375_),
    .B(_00478_),
    .C(_00479_),
    .Y(_00481_));
 sky130_fd_sc_hd__a21oi_1 _06646_ (.A1(_00478_),
    .A2(_00479_),
    .B1(_00375_),
    .Y(_00482_));
 sky130_fd_sc_hd__a211oi_2 _06647_ (.A1(_00359_),
    .A2(_00361_),
    .B1(_00480_),
    .C1(_00482_),
    .Y(_00483_));
 sky130_fd_sc_hd__o211a_1 _06648_ (.A1(_00480_),
    .A2(_00482_),
    .B1(_00359_),
    .C1(_00361_),
    .X(_00485_));
 sky130_fd_sc_hd__nor3_1 _06649_ (.A(_00256_),
    .B(_00483_),
    .C(_00485_),
    .Y(_00486_));
 sky130_fd_sc_hd__o21a_1 _06650_ (.A1(_00483_),
    .A2(_00485_),
    .B1(_00256_),
    .X(_00487_));
 sky130_fd_sc_hd__or2_1 _06651_ (.A(_00486_),
    .B(_00487_),
    .X(_00488_));
 sky130_fd_sc_hd__nor2_1 _06652_ (.A(_00363_),
    .B(_00488_),
    .Y(_00489_));
 sky130_fd_sc_hd__xor2_1 _06653_ (.A(_00363_),
    .B(_00488_),
    .X(_00490_));
 sky130_fd_sc_hd__and4bb_1 _06654_ (.A_N(_00243_),
    .B_N(_00488_),
    .C(_00365_),
    .D(_00363_),
    .X(_00491_));
 sky130_fd_sc_hd__xnor2_1 _06655_ (.A(_00367_),
    .B(_00490_),
    .Y(_00492_));
 sky130_fd_sc_hd__o21a_1 _06656_ (.A1(_00245_),
    .A2(_00247_),
    .B1(_00368_),
    .X(_00493_));
 sky130_fd_sc_hd__a21oi_1 _06657_ (.A1(_00255_),
    .A2(_00369_),
    .B1(_00493_),
    .Y(_00494_));
 sky130_fd_sc_hd__xor2_1 _06658_ (.A(_00492_),
    .B(_00494_),
    .X(net79));
 sky130_fd_sc_hd__or2_1 _06659_ (.A(_00405_),
    .B(_00408_),
    .X(_00496_));
 sky130_fd_sc_hd__or2_1 _06660_ (.A(_00377_),
    .B(_00384_),
    .X(_00497_));
 sky130_fd_sc_hd__nand3_1 _06661_ (.A(_00377_),
    .B(_00384_),
    .C(_00387_),
    .Y(_00498_));
 sky130_fd_sc_hd__and2_1 _06662_ (.A(_00497_),
    .B(_00498_),
    .X(_00499_));
 sky130_fd_sc_hd__and2_1 _06663_ (.A(_00496_),
    .B(_00499_),
    .X(_00500_));
 sky130_fd_sc_hd__xnor2_1 _06664_ (.A(_00496_),
    .B(_00499_),
    .Y(_00501_));
 sky130_fd_sc_hd__and4_1 _06665_ (.A(net518),
    .B(net605),
    .C(net333),
    .D(net325),
    .X(_00502_));
 sky130_fd_sc_hd__a22o_1 _06666_ (.A1(net519),
    .A2(net333),
    .B1(net325),
    .B2(net605),
    .X(_00503_));
 sky130_fd_sc_hd__and2b_1 _06667_ (.A_N(_00502_),
    .B(_00503_),
    .X(_00504_));
 sky130_fd_sc_hd__nand2_1 _06668_ (.A(net630),
    .B(net318),
    .Y(_00506_));
 sky130_fd_sc_hd__xnor2_1 _06669_ (.A(_00504_),
    .B(_00506_),
    .Y(_00507_));
 sky130_fd_sc_hd__and4_1 _06670_ (.A(net483),
    .B(net490),
    .C(net363),
    .D(net355),
    .X(_00508_));
 sky130_fd_sc_hd__a22o_1 _06671_ (.A1(net484),
    .A2(net364),
    .B1(net356),
    .B2(net490),
    .X(_00509_));
 sky130_fd_sc_hd__and2b_1 _06672_ (.A_N(_00508_),
    .B(_00509_),
    .X(_00510_));
 sky130_fd_sc_hd__nand2_1 _06673_ (.A(net499),
    .B(net338),
    .Y(_00511_));
 sky130_fd_sc_hd__xnor2_1 _06674_ (.A(_00510_),
    .B(_00511_),
    .Y(_00512_));
 sky130_fd_sc_hd__a31o_1 _06675_ (.A1(net519),
    .A2(net338),
    .A3(_00379_),
    .B1(_00378_),
    .X(_00513_));
 sky130_fd_sc_hd__and2_1 _06676_ (.A(_00512_),
    .B(_00513_),
    .X(_00514_));
 sky130_fd_sc_hd__xor2_1 _06677_ (.A(_00512_),
    .B(_00513_),
    .X(_00515_));
 sky130_fd_sc_hd__and2_1 _06678_ (.A(_00507_),
    .B(_00515_),
    .X(_00517_));
 sky130_fd_sc_hd__nor2_1 _06679_ (.A(_00507_),
    .B(_00515_),
    .Y(_00518_));
 sky130_fd_sc_hd__or2_1 _06680_ (.A(_00517_),
    .B(_00518_),
    .X(_00519_));
 sky130_fd_sc_hd__a31o_1 _06681_ (.A1(net483),
    .A2(net371),
    .A3(_00393_),
    .B1(_00391_),
    .X(_00520_));
 sky130_fd_sc_hd__o21bai_1 _06682_ (.A1(_00411_),
    .A2(_00413_),
    .B1_N(_00410_),
    .Y(_00521_));
 sky130_fd_sc_hd__nand4_1 _06683_ (.A(net460),
    .B(net453),
    .C(net394),
    .D(net378),
    .Y(_00522_));
 sky130_fd_sc_hd__a22o_1 _06684_ (.A1(net453),
    .A2(net394),
    .B1(net378),
    .B2(net460),
    .X(_00523_));
 sky130_fd_sc_hd__nand2_1 _06685_ (.A(net475),
    .B(net370),
    .Y(_00524_));
 sky130_fd_sc_hd__nand3b_1 _06686_ (.A_N(_00524_),
    .B(_00523_),
    .C(_00522_),
    .Y(_00525_));
 sky130_fd_sc_hd__a21bo_1 _06687_ (.A1(_00522_),
    .A2(_00523_),
    .B1_N(_00524_),
    .X(_00526_));
 sky130_fd_sc_hd__nand3_1 _06688_ (.A(_00521_),
    .B(_00525_),
    .C(_00526_),
    .Y(_00528_));
 sky130_fd_sc_hd__a21o_1 _06689_ (.A1(_00525_),
    .A2(_00526_),
    .B1(_00521_),
    .X(_00529_));
 sky130_fd_sc_hd__and3_1 _06690_ (.A(_00520_),
    .B(_00528_),
    .C(_00529_),
    .X(_00530_));
 sky130_fd_sc_hd__a21oi_1 _06691_ (.A1(_00528_),
    .A2(_00529_),
    .B1(_00520_),
    .Y(_00531_));
 sky130_fd_sc_hd__or2_1 _06692_ (.A(_00530_),
    .B(_00531_),
    .X(_00532_));
 sky130_fd_sc_hd__a21oi_2 _06693_ (.A1(_00397_),
    .A2(_00399_),
    .B1(_00532_),
    .Y(_00533_));
 sky130_fd_sc_hd__inv_2 _06694_ (.A(_00533_),
    .Y(_00534_));
 sky130_fd_sc_hd__and3_1 _06695_ (.A(_00397_),
    .B(_00399_),
    .C(_00532_),
    .X(_00535_));
 sky130_fd_sc_hd__nor3_1 _06696_ (.A(_00519_),
    .B(_00533_),
    .C(_00535_),
    .Y(_00536_));
 sky130_fd_sc_hd__or3_1 _06697_ (.A(_00519_),
    .B(_00533_),
    .C(_00535_),
    .X(_00537_));
 sky130_fd_sc_hd__o21a_1 _06698_ (.A1(_00533_),
    .A2(_00535_),
    .B1(_00519_),
    .X(_00539_));
 sky130_fd_sc_hd__a211oi_1 _06699_ (.A1(_00426_),
    .A2(_00430_),
    .B1(_00536_),
    .C1(_00539_),
    .Y(_00540_));
 sky130_fd_sc_hd__o211a_1 _06700_ (.A1(_00536_),
    .A2(_00539_),
    .B1(_00426_),
    .C1(_00430_),
    .X(_00541_));
 sky130_fd_sc_hd__a211oi_1 _06701_ (.A1(_00401_),
    .A2(_00403_),
    .B1(_00540_),
    .C1(_00541_),
    .Y(_00542_));
 sky130_fd_sc_hd__o211a_1 _06702_ (.A1(_00540_),
    .A2(_00541_),
    .B1(_00401_),
    .C1(_00403_),
    .X(_00543_));
 sky130_fd_sc_hd__a21o_1 _06703_ (.A1(_00432_),
    .A2(_00441_),
    .B1(_00439_),
    .X(_00544_));
 sky130_fd_sc_hd__and4_1 _06704_ (.A(net548),
    .B(net467),
    .C(net417),
    .D(net409),
    .X(_00545_));
 sky130_fd_sc_hd__a22o_1 _06705_ (.A1(net467),
    .A2(net417),
    .B1(net409),
    .B2(net548),
    .X(_00546_));
 sky130_fd_sc_hd__and2b_1 _06706_ (.A_N(_00545_),
    .B(_00546_),
    .X(_00547_));
 sky130_fd_sc_hd__nand2_1 _06707_ (.A(net447),
    .B(net402),
    .Y(_00548_));
 sky130_fd_sc_hd__xnor2_1 _06708_ (.A(_00547_),
    .B(_00548_),
    .Y(_00550_));
 sky130_fd_sc_hd__and4_1 _06709_ (.A(net190),
    .B(net432),
    .C(net300),
    .D(net224),
    .X(_00551_));
 sky130_fd_sc_hd__a22oi_2 _06710_ (.A1(net432),
    .A2(net300),
    .B1(net224),
    .B2(net190),
    .Y(_00552_));
 sky130_fd_sc_hd__nand2_1 _06711_ (.A(net424),
    .B(net387),
    .Y(_00553_));
 sky130_fd_sc_hd__or3_1 _06712_ (.A(_00551_),
    .B(_00552_),
    .C(_00553_),
    .X(_00554_));
 sky130_fd_sc_hd__o21ai_1 _06713_ (.A1(_00551_),
    .A2(_00552_),
    .B1(_00553_),
    .Y(_00555_));
 sky130_fd_sc_hd__a31o_1 _06714_ (.A1(net468),
    .A2(net424),
    .A3(_00416_),
    .B1(_00415_),
    .X(_00556_));
 sky130_fd_sc_hd__nand3_2 _06715_ (.A(_00554_),
    .B(_00555_),
    .C(_00556_),
    .Y(_00557_));
 sky130_fd_sc_hd__a21o_1 _06716_ (.A1(_00554_),
    .A2(_00555_),
    .B1(_00556_),
    .X(_00558_));
 sky130_fd_sc_hd__nand3_2 _06717_ (.A(_00550_),
    .B(_00557_),
    .C(_00558_),
    .Y(_00559_));
 sky130_fd_sc_hd__a21o_1 _06718_ (.A1(_00557_),
    .A2(_00558_),
    .B1(_00550_),
    .X(_00561_));
 sky130_fd_sc_hd__nand3_2 _06719_ (.A(_00544_),
    .B(_00559_),
    .C(_00561_),
    .Y(_00562_));
 sky130_fd_sc_hd__a21o_1 _06720_ (.A1(_00559_),
    .A2(_00561_),
    .B1(_00544_),
    .X(_00563_));
 sky130_fd_sc_hd__o211ai_2 _06721_ (.A1(_00422_),
    .A2(_00424_),
    .B1(_00562_),
    .C1(_00563_),
    .Y(_00564_));
 sky130_fd_sc_hd__a211o_1 _06722_ (.A1(_00562_),
    .A2(_00563_),
    .B1(_00422_),
    .C1(_00424_),
    .X(_00565_));
 sky130_fd_sc_hd__nand2_1 _06723_ (.A(_00564_),
    .B(_00565_),
    .Y(_00566_));
 sky130_fd_sc_hd__nand2_1 _06724_ (.A(_00434_),
    .B(_00437_),
    .Y(_00567_));
 sky130_fd_sc_hd__o21bai_1 _06725_ (.A1(_00444_),
    .A2(_00446_),
    .B1_N(_00445_),
    .Y(_00568_));
 sky130_fd_sc_hd__and4_1 _06726_ (.A(net212),
    .B(net203),
    .C(net172),
    .D(net164),
    .X(_00569_));
 sky130_fd_sc_hd__a22oi_1 _06727_ (.A1(net203),
    .A2(net172),
    .B1(net164),
    .B2(net212),
    .Y(_00570_));
 sky130_fd_sc_hd__nand2_1 _06728_ (.A(net195),
    .B(net179),
    .Y(_00572_));
 sky130_fd_sc_hd__or3_1 _06729_ (.A(_00569_),
    .B(_00570_),
    .C(_00572_),
    .X(_00573_));
 sky130_fd_sc_hd__o21ai_1 _06730_ (.A1(_00569_),
    .A2(_00570_),
    .B1(_00572_),
    .Y(_00574_));
 sky130_fd_sc_hd__and3_1 _06731_ (.A(_00568_),
    .B(_00573_),
    .C(_00574_),
    .X(_00575_));
 sky130_fd_sc_hd__a21o_1 _06732_ (.A1(_00573_),
    .A2(_00574_),
    .B1(_00568_),
    .X(_00576_));
 sky130_fd_sc_hd__and2b_1 _06733_ (.A_N(_00575_),
    .B(_00576_),
    .X(_00577_));
 sky130_fd_sc_hd__xor2_1 _06734_ (.A(_00567_),
    .B(_00577_),
    .X(_00578_));
 sky130_fd_sc_hd__nand2_1 _06735_ (.A(net218),
    .B(net621),
    .Y(_00579_));
 sky130_fd_sc_hd__and4_1 _06736_ (.A(net240),
    .B(net233),
    .C(net613),
    .D(net596),
    .X(_00580_));
 sky130_fd_sc_hd__a22oi_1 _06737_ (.A1(net233),
    .A2(net613),
    .B1(net596),
    .B2(net240),
    .Y(_00581_));
 sky130_fd_sc_hd__nor2_1 _06738_ (.A(_00580_),
    .B(_00581_),
    .Y(_00583_));
 sky130_fd_sc_hd__xnor2_1 _06739_ (.A(_00579_),
    .B(_00583_),
    .Y(_00584_));
 sky130_fd_sc_hd__nand2_1 _06740_ (.A(net258),
    .B(net590),
    .Y(_00585_));
 sky130_fd_sc_hd__and4_1 _06741_ (.A(net437),
    .B(net345),
    .C(net581),
    .D(net575),
    .X(_00586_));
 sky130_fd_sc_hd__a22oi_2 _06742_ (.A1(net348),
    .A2(net581),
    .B1(net575),
    .B2(net437),
    .Y(_00587_));
 sky130_fd_sc_hd__or3_1 _06743_ (.A(_00585_),
    .B(_00586_),
    .C(_00587_),
    .X(_00588_));
 sky130_fd_sc_hd__o21ai_1 _06744_ (.A1(_00586_),
    .A2(_00587_),
    .B1(_00585_),
    .Y(_00589_));
 sky130_fd_sc_hd__o21bai_1 _06745_ (.A1(_00449_),
    .A2(_00452_),
    .B1_N(_00450_),
    .Y(_00590_));
 sky130_fd_sc_hd__nand3_1 _06746_ (.A(_00588_),
    .B(_00589_),
    .C(_00590_),
    .Y(_00591_));
 sky130_fd_sc_hd__a21o_1 _06747_ (.A1(_00588_),
    .A2(_00589_),
    .B1(_00590_),
    .X(_00592_));
 sky130_fd_sc_hd__nand3_1 _06748_ (.A(_00584_),
    .B(_00591_),
    .C(_00592_),
    .Y(_00594_));
 sky130_fd_sc_hd__a21o_1 _06749_ (.A1(_00591_),
    .A2(_00592_),
    .B1(_00584_),
    .X(_00595_));
 sky130_fd_sc_hd__a21bo_1 _06750_ (.A1(_00448_),
    .A2(_00457_),
    .B1_N(_00456_),
    .X(_00596_));
 sky130_fd_sc_hd__nand3_2 _06751_ (.A(_00594_),
    .B(_00595_),
    .C(_00596_),
    .Y(_00597_));
 sky130_fd_sc_hd__a21o_1 _06752_ (.A1(_00594_),
    .A2(_00595_),
    .B1(_00596_),
    .X(_00598_));
 sky130_fd_sc_hd__and3_1 _06753_ (.A(_00578_),
    .B(_00597_),
    .C(_00598_),
    .X(_00599_));
 sky130_fd_sc_hd__nand3_1 _06754_ (.A(_00578_),
    .B(_00597_),
    .C(_00598_),
    .Y(_00600_));
 sky130_fd_sc_hd__a21oi_2 _06755_ (.A1(_00597_),
    .A2(_00598_),
    .B1(_00578_),
    .Y(_00601_));
 sky130_fd_sc_hd__a211oi_4 _06756_ (.A1(_00461_),
    .A2(_00465_),
    .B1(_00599_),
    .C1(_00601_),
    .Y(_00602_));
 sky130_fd_sc_hd__o211a_1 _06757_ (.A1(_00599_),
    .A2(_00601_),
    .B1(_00461_),
    .C1(_00465_),
    .X(_00603_));
 sky130_fd_sc_hd__nor3_1 _06758_ (.A(_00566_),
    .B(_00602_),
    .C(_00603_),
    .Y(_00605_));
 sky130_fd_sc_hd__or3_2 _06759_ (.A(_00566_),
    .B(_00602_),
    .C(_00603_),
    .X(_00606_));
 sky130_fd_sc_hd__o21ai_2 _06760_ (.A1(_00602_),
    .A2(_00603_),
    .B1(_00566_),
    .Y(_00607_));
 sky130_fd_sc_hd__o211ai_4 _06761_ (.A1(_00467_),
    .A2(net147),
    .B1(_00606_),
    .C1(_00607_),
    .Y(_00608_));
 sky130_fd_sc_hd__a211o_1 _06762_ (.A1(_00606_),
    .A2(_00607_),
    .B1(_00467_),
    .C1(_00469_),
    .X(_00609_));
 sky130_fd_sc_hd__and4bb_1 _06763_ (.A_N(_00542_),
    .B_N(_00543_),
    .C(_00608_),
    .D(_00609_),
    .X(_00610_));
 sky130_fd_sc_hd__or4bb_1 _06764_ (.A(_00542_),
    .B(_00543_),
    .C_N(_00608_),
    .D_N(_00609_),
    .X(_00611_));
 sky130_fd_sc_hd__a2bb2oi_1 _06765_ (.A1_N(_00542_),
    .A2_N(_00543_),
    .B1(_00608_),
    .B2(_00609_),
    .Y(_00612_));
 sky130_fd_sc_hd__a211oi_2 _06766_ (.A1(_00472_),
    .A2(_00476_),
    .B1(_00610_),
    .C1(_00612_),
    .Y(_00613_));
 sky130_fd_sc_hd__o211a_1 _06767_ (.A1(_00610_),
    .A2(_00612_),
    .B1(_00472_),
    .C1(_00476_),
    .X(_00614_));
 sky130_fd_sc_hd__nor3_2 _06768_ (.A(_00501_),
    .B(_00613_),
    .C(_00614_),
    .Y(_00616_));
 sky130_fd_sc_hd__o21a_1 _06769_ (.A1(_00613_),
    .A2(_00614_),
    .B1(_00501_),
    .X(_00617_));
 sky130_fd_sc_hd__a211oi_1 _06770_ (.A1(_00478_),
    .A2(_00481_),
    .B1(_00616_),
    .C1(_00617_),
    .Y(_00618_));
 sky130_fd_sc_hd__a211o_1 _06771_ (.A1(_00478_),
    .A2(_00481_),
    .B1(_00616_),
    .C1(_00617_),
    .X(_00619_));
 sky130_fd_sc_hd__o211ai_1 _06772_ (.A1(_00616_),
    .A2(_00617_),
    .B1(_00478_),
    .C1(_00481_),
    .Y(_00620_));
 sky130_fd_sc_hd__and3_1 _06773_ (.A(_00372_),
    .B(_00619_),
    .C(_00620_),
    .X(_00621_));
 sky130_fd_sc_hd__nand3_1 _06774_ (.A(_00372_),
    .B(_00619_),
    .C(_00620_),
    .Y(_00622_));
 sky130_fd_sc_hd__a21o_1 _06775_ (.A1(_00619_),
    .A2(_00620_),
    .B1(_00372_),
    .X(_00623_));
 sky130_fd_sc_hd__o211ai_2 _06776_ (.A1(_00483_),
    .A2(_00486_),
    .B1(_00622_),
    .C1(_00623_),
    .Y(_00624_));
 sky130_fd_sc_hd__a211o_1 _06777_ (.A1(_00622_),
    .A2(_00623_),
    .B1(_00483_),
    .C1(_00486_),
    .X(_00625_));
 sky130_fd_sc_hd__and2_1 _06778_ (.A(_00624_),
    .B(_00625_),
    .X(_00627_));
 sky130_fd_sc_hd__xor2_1 _06779_ (.A(_00489_),
    .B(_00627_),
    .X(_00628_));
 sky130_fd_sc_hd__o21ba_1 _06780_ (.A1(_00492_),
    .A2(_00494_),
    .B1_N(_00491_),
    .X(_00629_));
 sky130_fd_sc_hd__xnor2_1 _06781_ (.A(_00628_),
    .B(_00629_),
    .Y(net80));
 sky130_fd_sc_hd__or2_1 _06782_ (.A(_00540_),
    .B(_00542_),
    .X(_00630_));
 sky130_fd_sc_hd__a31o_1 _06783_ (.A1(net630),
    .A2(net318),
    .A3(_00503_),
    .B1(_00502_),
    .X(_00631_));
 sky130_fd_sc_hd__and3_1 _06784_ (.A(net630),
    .B(net310),
    .C(_00631_),
    .X(_00632_));
 sky130_fd_sc_hd__a21oi_1 _06785_ (.A1(net630),
    .A2(net310),
    .B1(_00631_),
    .Y(_00633_));
 sky130_fd_sc_hd__nor2_1 _06786_ (.A(_00632_),
    .B(_00633_),
    .Y(_00634_));
 sky130_fd_sc_hd__o21ai_1 _06787_ (.A1(_00514_),
    .A2(_00517_),
    .B1(_00634_),
    .Y(_00635_));
 sky130_fd_sc_hd__or3_1 _06788_ (.A(_00514_),
    .B(_00517_),
    .C(_00634_),
    .X(_00637_));
 sky130_fd_sc_hd__and2_1 _06789_ (.A(_00635_),
    .B(_00637_),
    .X(_00638_));
 sky130_fd_sc_hd__and2b_1 _06790_ (.A_N(_00497_),
    .B(_00638_),
    .X(_00639_));
 sky130_fd_sc_hd__xnor2_1 _06791_ (.A(_00497_),
    .B(_00638_),
    .Y(_00640_));
 sky130_fd_sc_hd__nand2_1 _06792_ (.A(_00630_),
    .B(_00640_),
    .Y(_00641_));
 sky130_fd_sc_hd__xnor2_1 _06793_ (.A(_00630_),
    .B(_00640_),
    .Y(_00642_));
 sky130_fd_sc_hd__and4_1 _06794_ (.A(net498),
    .B(net518),
    .C(net332),
    .D(net326),
    .X(_00643_));
 sky130_fd_sc_hd__a22oi_1 _06795_ (.A1(net498),
    .A2(net332),
    .B1(net326),
    .B2(net518),
    .Y(_00644_));
 sky130_fd_sc_hd__nor2_1 _06796_ (.A(_00643_),
    .B(_00644_),
    .Y(_00645_));
 sky130_fd_sc_hd__nand2_1 _06797_ (.A(net605),
    .B(net318),
    .Y(_00646_));
 sky130_fd_sc_hd__xnor2_1 _06798_ (.A(_00645_),
    .B(_00646_),
    .Y(_00648_));
 sky130_fd_sc_hd__and4_1 _06799_ (.A(net484),
    .B(net476),
    .C(net363),
    .D(net355),
    .X(_00649_));
 sky130_fd_sc_hd__a22oi_2 _06800_ (.A1(net476),
    .A2(net364),
    .B1(net356),
    .B2(net484),
    .Y(_00650_));
 sky130_fd_sc_hd__nand2_1 _06801_ (.A(net491),
    .B(net338),
    .Y(_00651_));
 sky130_fd_sc_hd__or3_1 _06802_ (.A(_00649_),
    .B(_00650_),
    .C(_00651_),
    .X(_00652_));
 sky130_fd_sc_hd__o21ai_1 _06803_ (.A1(_00649_),
    .A2(_00650_),
    .B1(_00651_),
    .Y(_00653_));
 sky130_fd_sc_hd__a31o_1 _06804_ (.A1(net499),
    .A2(net338),
    .A3(_00509_),
    .B1(_00508_),
    .X(_00654_));
 sky130_fd_sc_hd__and3_1 _06805_ (.A(_00652_),
    .B(_00653_),
    .C(_00654_),
    .X(_00655_));
 sky130_fd_sc_hd__a21oi_1 _06806_ (.A1(_00652_),
    .A2(_00653_),
    .B1(_00654_),
    .Y(_00656_));
 sky130_fd_sc_hd__nor3b_1 _06807_ (.A(_00655_),
    .B(_00656_),
    .C_N(_00648_),
    .Y(_00657_));
 sky130_fd_sc_hd__o21ba_1 _06808_ (.A1(_00655_),
    .A2(_00656_),
    .B1_N(_00648_),
    .X(_00659_));
 sky130_fd_sc_hd__or2_1 _06809_ (.A(_00657_),
    .B(_00659_),
    .X(_00660_));
 sky130_fd_sc_hd__nand2_1 _06810_ (.A(_00522_),
    .B(_00525_),
    .Y(_00661_));
 sky130_fd_sc_hd__a31o_1 _06811_ (.A1(net447),
    .A2(net402),
    .A3(_00546_),
    .B1(_00545_),
    .X(_00662_));
 sky130_fd_sc_hd__nand4_1 _06812_ (.A(net453),
    .B(net447),
    .C(net394),
    .D(net378),
    .Y(_00663_));
 sky130_fd_sc_hd__a22o_1 _06813_ (.A1(net447),
    .A2(net394),
    .B1(net378),
    .B2(net453),
    .X(_00664_));
 sky130_fd_sc_hd__nand2_1 _06814_ (.A(net460),
    .B(net370),
    .Y(_00665_));
 sky130_fd_sc_hd__nand3b_1 _06815_ (.A_N(_00665_),
    .B(_00664_),
    .C(_00663_),
    .Y(_00666_));
 sky130_fd_sc_hd__a21bo_1 _06816_ (.A1(_00663_),
    .A2(_00664_),
    .B1_N(_00665_),
    .X(_00667_));
 sky130_fd_sc_hd__nand3_1 _06817_ (.A(_00662_),
    .B(_00666_),
    .C(_00667_),
    .Y(_00668_));
 sky130_fd_sc_hd__a21o_1 _06818_ (.A1(_00666_),
    .A2(_00667_),
    .B1(_00662_),
    .X(_00670_));
 sky130_fd_sc_hd__nand3_1 _06819_ (.A(_00661_),
    .B(_00668_),
    .C(_00670_),
    .Y(_00671_));
 sky130_fd_sc_hd__a21o_1 _06820_ (.A1(_00668_),
    .A2(_00670_),
    .B1(_00661_),
    .X(_00672_));
 sky130_fd_sc_hd__a21bo_1 _06821_ (.A1(_00520_),
    .A2(_00529_),
    .B1_N(_00528_),
    .X(_00673_));
 sky130_fd_sc_hd__and3_1 _06822_ (.A(_00671_),
    .B(_00672_),
    .C(_00673_),
    .X(_00674_));
 sky130_fd_sc_hd__inv_2 _06823_ (.A(_00674_),
    .Y(_00675_));
 sky130_fd_sc_hd__a21oi_1 _06824_ (.A1(_00671_),
    .A2(_00672_),
    .B1(_00673_),
    .Y(_00676_));
 sky130_fd_sc_hd__nor3_1 _06825_ (.A(_00660_),
    .B(_00674_),
    .C(_00676_),
    .Y(_00677_));
 sky130_fd_sc_hd__or3_1 _06826_ (.A(_00660_),
    .B(_00674_),
    .C(_00676_),
    .X(_00678_));
 sky130_fd_sc_hd__o21a_1 _06827_ (.A1(_00674_),
    .A2(_00676_),
    .B1(_00660_),
    .X(_00679_));
 sky130_fd_sc_hd__a211oi_2 _06828_ (.A1(_00562_),
    .A2(_00564_),
    .B1(_00677_),
    .C1(_00679_),
    .Y(_00681_));
 sky130_fd_sc_hd__o211a_1 _06829_ (.A1(_00677_),
    .A2(_00679_),
    .B1(_00562_),
    .C1(_00564_),
    .X(_00682_));
 sky130_fd_sc_hd__a211oi_2 _06830_ (.A1(_00534_),
    .A2(_00537_),
    .B1(_00681_),
    .C1(_00682_),
    .Y(_00683_));
 sky130_fd_sc_hd__o211a_1 _06831_ (.A1(_00681_),
    .A2(_00682_),
    .B1(_00534_),
    .C1(_00537_),
    .X(_00684_));
 sky130_fd_sc_hd__a21o_1 _06832_ (.A1(_00567_),
    .A2(_00576_),
    .B1(_00575_),
    .X(_00685_));
 sky130_fd_sc_hd__and4_1 _06833_ (.A(net467),
    .B(net387),
    .C(net417),
    .D(net409),
    .X(_00686_));
 sky130_fd_sc_hd__a22o_1 _06834_ (.A1(net387),
    .A2(net417),
    .B1(net409),
    .B2(net467),
    .X(_00687_));
 sky130_fd_sc_hd__and2b_1 _06835_ (.A_N(_00686_),
    .B(_00687_),
    .X(_00688_));
 sky130_fd_sc_hd__nand2_1 _06836_ (.A(net548),
    .B(net402),
    .Y(_00689_));
 sky130_fd_sc_hd__xnor2_1 _06837_ (.A(_00688_),
    .B(_00689_),
    .Y(_00690_));
 sky130_fd_sc_hd__nand4_1 _06838_ (.A(net190),
    .B(net432),
    .C(net224),
    .D(net181),
    .Y(_00692_));
 sky130_fd_sc_hd__a22o_1 _06839_ (.A1(net432),
    .A2(net224),
    .B1(net181),
    .B2(net190),
    .X(_00693_));
 sky130_fd_sc_hd__nand2_1 _06840_ (.A(net424),
    .B(net303),
    .Y(_00694_));
 sky130_fd_sc_hd__nand3b_1 _06841_ (.A_N(_00694_),
    .B(_00693_),
    .C(_00692_),
    .Y(_00695_));
 sky130_fd_sc_hd__a21bo_1 _06842_ (.A1(_00692_),
    .A2(_00693_),
    .B1_N(_00694_),
    .X(_00696_));
 sky130_fd_sc_hd__o21bai_1 _06843_ (.A1(_00552_),
    .A2(_00553_),
    .B1_N(_00551_),
    .Y(_00697_));
 sky130_fd_sc_hd__nand3_2 _06844_ (.A(_00695_),
    .B(_00696_),
    .C(_00697_),
    .Y(_00698_));
 sky130_fd_sc_hd__a21o_1 _06845_ (.A1(_00695_),
    .A2(_00696_),
    .B1(_00697_),
    .X(_00699_));
 sky130_fd_sc_hd__nand3_2 _06846_ (.A(_00690_),
    .B(_00698_),
    .C(_00699_),
    .Y(_00700_));
 sky130_fd_sc_hd__a21o_1 _06847_ (.A1(_00698_),
    .A2(_00699_),
    .B1(_00690_),
    .X(_00701_));
 sky130_fd_sc_hd__and3_1 _06848_ (.A(_00685_),
    .B(_00700_),
    .C(_00701_),
    .X(_00703_));
 sky130_fd_sc_hd__a21oi_1 _06849_ (.A1(_00700_),
    .A2(_00701_),
    .B1(_00685_),
    .Y(_00704_));
 sky130_fd_sc_hd__a211oi_2 _06850_ (.A1(_00557_),
    .A2(_00559_),
    .B1(_00703_),
    .C1(_00704_),
    .Y(_00705_));
 sky130_fd_sc_hd__o211a_1 _06851_ (.A1(_00703_),
    .A2(_00704_),
    .B1(_00557_),
    .C1(_00559_),
    .X(_00706_));
 sky130_fd_sc_hd__and2b_1 _06852_ (.A_N(_00569_),
    .B(_00573_),
    .X(_00707_));
 sky130_fd_sc_hd__o21ba_1 _06853_ (.A1(_00579_),
    .A2(_00581_),
    .B1_N(_00580_),
    .X(_00708_));
 sky130_fd_sc_hd__and4_1 _06854_ (.A(net212),
    .B(net203),
    .C(net164),
    .D(net621),
    .X(_00709_));
 sky130_fd_sc_hd__a22oi_1 _06855_ (.A1(net203),
    .A2(net164),
    .B1(net621),
    .B2(net212),
    .Y(_00710_));
 sky130_fd_sc_hd__nor2_1 _06856_ (.A(_00709_),
    .B(_00710_),
    .Y(_00711_));
 sky130_fd_sc_hd__nand2_1 _06857_ (.A(net195),
    .B(net172),
    .Y(_00712_));
 sky130_fd_sc_hd__xnor2_1 _06858_ (.A(_00711_),
    .B(_00712_),
    .Y(_00714_));
 sky130_fd_sc_hd__nand2b_1 _06859_ (.A_N(_00708_),
    .B(_00714_),
    .Y(_00715_));
 sky130_fd_sc_hd__xnor2_1 _06860_ (.A(_00708_),
    .B(_00714_),
    .Y(_00716_));
 sky130_fd_sc_hd__nand2b_1 _06861_ (.A_N(_00707_),
    .B(_00716_),
    .Y(_00717_));
 sky130_fd_sc_hd__xnor2_1 _06862_ (.A(_00707_),
    .B(_00716_),
    .Y(_00718_));
 sky130_fd_sc_hd__and4_1 _06863_ (.A(net240),
    .B(net233),
    .C(net597),
    .D(net590),
    .X(_00719_));
 sky130_fd_sc_hd__a22oi_1 _06864_ (.A1(net233),
    .A2(net597),
    .B1(net590),
    .B2(net240),
    .Y(_00720_));
 sky130_fd_sc_hd__nor2_1 _06865_ (.A(_00719_),
    .B(_00720_),
    .Y(_00721_));
 sky130_fd_sc_hd__nand2_1 _06866_ (.A(net218),
    .B(net613),
    .Y(_00722_));
 sky130_fd_sc_hd__xnor2_1 _06867_ (.A(_00721_),
    .B(_00722_),
    .Y(_00723_));
 sky130_fd_sc_hd__nand2_1 _06868_ (.A(net258),
    .B(net582),
    .Y(_00725_));
 sky130_fd_sc_hd__and4_1 _06869_ (.A(net437),
    .B(net345),
    .C(net16),
    .D(net568),
    .X(_00726_));
 sky130_fd_sc_hd__a22oi_2 _06870_ (.A1(net345),
    .A2(net576),
    .B1(net568),
    .B2(net437),
    .Y(_00727_));
 sky130_fd_sc_hd__or3_1 _06871_ (.A(_00725_),
    .B(_00726_),
    .C(_00727_),
    .X(_00728_));
 sky130_fd_sc_hd__o21ai_1 _06872_ (.A1(_00726_),
    .A2(_00727_),
    .B1(_00725_),
    .Y(_00729_));
 sky130_fd_sc_hd__o21bai_1 _06873_ (.A1(_00585_),
    .A2(_00587_),
    .B1_N(_00586_),
    .Y(_00730_));
 sky130_fd_sc_hd__nand3_1 _06874_ (.A(_00728_),
    .B(_00729_),
    .C(_00730_),
    .Y(_00731_));
 sky130_fd_sc_hd__a21o_1 _06875_ (.A1(_00728_),
    .A2(_00729_),
    .B1(_00730_),
    .X(_00732_));
 sky130_fd_sc_hd__nand3_1 _06876_ (.A(_00723_),
    .B(_00731_),
    .C(_00732_),
    .Y(_00733_));
 sky130_fd_sc_hd__a21o_1 _06877_ (.A1(_00731_),
    .A2(_00732_),
    .B1(_00723_),
    .X(_00734_));
 sky130_fd_sc_hd__a21bo_1 _06878_ (.A1(_00584_),
    .A2(_00592_),
    .B1_N(_00591_),
    .X(_00736_));
 sky130_fd_sc_hd__nand3_2 _06879_ (.A(_00733_),
    .B(_00734_),
    .C(_00736_),
    .Y(_00737_));
 sky130_fd_sc_hd__a21o_1 _06880_ (.A1(_00733_),
    .A2(_00734_),
    .B1(_00736_),
    .X(_00738_));
 sky130_fd_sc_hd__and3_1 _06881_ (.A(_00718_),
    .B(_00737_),
    .C(_00738_),
    .X(_00739_));
 sky130_fd_sc_hd__nand3_1 _06882_ (.A(_00718_),
    .B(_00737_),
    .C(_00738_),
    .Y(_00740_));
 sky130_fd_sc_hd__a21oi_1 _06883_ (.A1(_00737_),
    .A2(_00738_),
    .B1(_00718_),
    .Y(_00741_));
 sky130_fd_sc_hd__a211o_1 _06884_ (.A1(_00597_),
    .A2(_00600_),
    .B1(_00739_),
    .C1(_00741_),
    .X(_00742_));
 sky130_fd_sc_hd__o211ai_1 _06885_ (.A1(_00739_),
    .A2(_00741_),
    .B1(_00597_),
    .C1(_00600_),
    .Y(_00743_));
 sky130_fd_sc_hd__or4bb_2 _06886_ (.A(_00705_),
    .B(_00706_),
    .C_N(_00742_),
    .D_N(_00743_),
    .X(_00744_));
 sky130_fd_sc_hd__a2bb2o_1 _06887_ (.A1_N(_00705_),
    .A2_N(_00706_),
    .B1(_00742_),
    .B2(_00743_),
    .X(_00745_));
 sky130_fd_sc_hd__o211a_1 _06888_ (.A1(_00602_),
    .A2(_00605_),
    .B1(_00744_),
    .C1(_00745_),
    .X(_00747_));
 sky130_fd_sc_hd__a211oi_1 _06889_ (.A1(_00744_),
    .A2(_00745_),
    .B1(_00602_),
    .C1(_00605_),
    .Y(_00748_));
 sky130_fd_sc_hd__nor4_1 _06890_ (.A(_00683_),
    .B(_00684_),
    .C(_00747_),
    .D(_00748_),
    .Y(_00749_));
 sky130_fd_sc_hd__o22a_1 _06891_ (.A1(_00683_),
    .A2(_00684_),
    .B1(_00747_),
    .B2(_00748_),
    .X(_00750_));
 sky130_fd_sc_hd__a211oi_2 _06892_ (.A1(_00608_),
    .A2(_00611_),
    .B1(net141),
    .C1(_00750_),
    .Y(_00751_));
 sky130_fd_sc_hd__o211a_1 _06893_ (.A1(net141),
    .A2(_00750_),
    .B1(_00608_),
    .C1(_00611_),
    .X(_00752_));
 sky130_fd_sc_hd__nor3_1 _06894_ (.A(_00642_),
    .B(_00751_),
    .C(_00752_),
    .Y(_00753_));
 sky130_fd_sc_hd__or3_1 _06895_ (.A(_00642_),
    .B(_00751_),
    .C(_00752_),
    .X(_00754_));
 sky130_fd_sc_hd__o21ai_1 _06896_ (.A1(_00751_),
    .A2(_00752_),
    .B1(_00642_),
    .Y(_00755_));
 sky130_fd_sc_hd__o211ai_2 _06897_ (.A1(_00613_),
    .A2(_00616_),
    .B1(_00754_),
    .C1(_00755_),
    .Y(_00756_));
 sky130_fd_sc_hd__a211o_1 _06898_ (.A1(_00754_),
    .A2(_00755_),
    .B1(_00613_),
    .C1(_00616_),
    .X(_00758_));
 sky130_fd_sc_hd__nand3_1 _06899_ (.A(_00500_),
    .B(_00756_),
    .C(_00758_),
    .Y(_00759_));
 sky130_fd_sc_hd__a21o_1 _06900_ (.A1(_00756_),
    .A2(_00758_),
    .B1(_00500_),
    .X(_00760_));
 sky130_fd_sc_hd__o211a_1 _06901_ (.A1(_00618_),
    .A2(_00621_),
    .B1(_00759_),
    .C1(_00760_),
    .X(_00761_));
 sky130_fd_sc_hd__a211o_1 _06902_ (.A1(_00759_),
    .A2(_00760_),
    .B1(_00618_),
    .C1(_00621_),
    .X(_00762_));
 sky130_fd_sc_hd__and2b_1 _06903_ (.A_N(_00761_),
    .B(_00762_),
    .X(_00763_));
 sky130_fd_sc_hd__and2b_1 _06904_ (.A_N(_00624_),
    .B(_00763_),
    .X(_00764_));
 sky130_fd_sc_hd__xor2_1 _06905_ (.A(_00624_),
    .B(_00763_),
    .X(_00765_));
 sky130_fd_sc_hd__and4bb_1 _06906_ (.A_N(_00249_),
    .B_N(_00492_),
    .C(_00628_),
    .D(_00369_),
    .X(_00766_));
 sky130_fd_sc_hd__o21ai_1 _06907_ (.A1(_00489_),
    .A2(_00491_),
    .B1(_00627_),
    .Y(_00767_));
 sky130_fd_sc_hd__inv_2 _06908_ (.A(_00767_),
    .Y(_00769_));
 sky130_fd_sc_hd__and3b_1 _06909_ (.A_N(_00492_),
    .B(_00493_),
    .C(_00628_),
    .X(_00770_));
 sky130_fd_sc_hd__a211o_1 _06910_ (.A1(_00252_),
    .A2(_00766_),
    .B1(_00769_),
    .C1(_00770_),
    .X(_00771_));
 sky130_fd_sc_hd__and3_1 _06911_ (.A(_00041_),
    .B(_00250_),
    .C(_00766_),
    .X(_00772_));
 sky130_fd_sc_hd__a21oi_2 _06912_ (.A1(_00253_),
    .A2(_00766_),
    .B1(_00771_),
    .Y(_00773_));
 sky130_fd_sc_hd__xor2_1 _06913_ (.A(_00765_),
    .B(_00773_),
    .X(net81));
 sky130_fd_sc_hd__nor2_1 _06914_ (.A(_00655_),
    .B(_00657_),
    .Y(_00774_));
 sky130_fd_sc_hd__a31o_1 _06915_ (.A1(net605),
    .A2(net318),
    .A3(_00645_),
    .B1(_00643_),
    .X(_00775_));
 sky130_fd_sc_hd__a22o_1 _06916_ (.A1(net605),
    .A2(net310),
    .B1(net296),
    .B2(net628),
    .X(_00776_));
 sky130_fd_sc_hd__and4_1 _06917_ (.A(net602),
    .B(net628),
    .C(net310),
    .D(net296),
    .X(_00777_));
 sky130_fd_sc_hd__inv_2 _06918_ (.A(_00777_),
    .Y(_00779_));
 sky130_fd_sc_hd__and3_1 _06919_ (.A(_00775_),
    .B(_00776_),
    .C(_00779_),
    .X(_00780_));
 sky130_fd_sc_hd__a21oi_1 _06920_ (.A1(_00776_),
    .A2(_00779_),
    .B1(_00775_),
    .Y(_00781_));
 sky130_fd_sc_hd__nor2_1 _06921_ (.A(_00780_),
    .B(_00781_),
    .Y(_00782_));
 sky130_fd_sc_hd__or3_1 _06922_ (.A(_00774_),
    .B(_00780_),
    .C(_00781_),
    .X(_00783_));
 sky130_fd_sc_hd__xnor2_1 _06923_ (.A(_00774_),
    .B(_00782_),
    .Y(_00784_));
 sky130_fd_sc_hd__nand2_1 _06924_ (.A(_00632_),
    .B(_00784_),
    .Y(_00785_));
 sky130_fd_sc_hd__xnor2_1 _06925_ (.A(_00632_),
    .B(_00784_),
    .Y(_00786_));
 sky130_fd_sc_hd__nor2_1 _06926_ (.A(_00635_),
    .B(_00786_),
    .Y(_00787_));
 sky130_fd_sc_hd__xor2_1 _06927_ (.A(_00635_),
    .B(_00786_),
    .X(_00788_));
 sky130_fd_sc_hd__nor3_1 _06928_ (.A(_00681_),
    .B(_00683_),
    .C(_00788_),
    .Y(_00790_));
 sky130_fd_sc_hd__o21a_1 _06929_ (.A1(_00681_),
    .A2(_00683_),
    .B1(_00788_),
    .X(_00791_));
 sky130_fd_sc_hd__nor2_1 _06930_ (.A(_00790_),
    .B(_00791_),
    .Y(_00792_));
 sky130_fd_sc_hd__and2_1 _06931_ (.A(_00639_),
    .B(_00792_),
    .X(_00793_));
 sky130_fd_sc_hd__xnor2_1 _06932_ (.A(_00639_),
    .B(_00792_),
    .Y(_00794_));
 sky130_fd_sc_hd__nand2_1 _06933_ (.A(net518),
    .B(net318),
    .Y(_00795_));
 sky130_fd_sc_hd__and4_1 _06934_ (.A(net490),
    .B(net498),
    .C(net332),
    .D(net325),
    .X(_00796_));
 sky130_fd_sc_hd__a22o_1 _06935_ (.A1(net490),
    .A2(net332),
    .B1(net325),
    .B2(net498),
    .X(_00797_));
 sky130_fd_sc_hd__and2b_1 _06936_ (.A_N(_00796_),
    .B(_00797_),
    .X(_00798_));
 sky130_fd_sc_hd__xnor2_1 _06937_ (.A(_00795_),
    .B(_00798_),
    .Y(_00799_));
 sky130_fd_sc_hd__nand2_1 _06938_ (.A(net484),
    .B(net338),
    .Y(_00801_));
 sky130_fd_sc_hd__and4_1 _06939_ (.A(net476),
    .B(net461),
    .C(net363),
    .D(net355),
    .X(_00802_));
 sky130_fd_sc_hd__a22oi_2 _06940_ (.A1(net461),
    .A2(net363),
    .B1(net355),
    .B2(net476),
    .Y(_00803_));
 sky130_fd_sc_hd__or3_1 _06941_ (.A(_00801_),
    .B(_00802_),
    .C(_00803_),
    .X(_00804_));
 sky130_fd_sc_hd__o21ai_1 _06942_ (.A1(_00802_),
    .A2(_00803_),
    .B1(_00801_),
    .Y(_00805_));
 sky130_fd_sc_hd__o21bai_1 _06943_ (.A1(_00650_),
    .A2(_00651_),
    .B1_N(_00649_),
    .Y(_00806_));
 sky130_fd_sc_hd__and3_1 _06944_ (.A(_00804_),
    .B(_00805_),
    .C(_00806_),
    .X(_00807_));
 sky130_fd_sc_hd__a21o_1 _06945_ (.A1(_00804_),
    .A2(_00805_),
    .B1(_00806_),
    .X(_00808_));
 sky130_fd_sc_hd__and2b_1 _06946_ (.A_N(_00807_),
    .B(_00808_),
    .X(_00809_));
 sky130_fd_sc_hd__xnor2_1 _06947_ (.A(_00799_),
    .B(_00809_),
    .Y(_00810_));
 sky130_fd_sc_hd__nand2_1 _06948_ (.A(_00663_),
    .B(_00666_),
    .Y(_00812_));
 sky130_fd_sc_hd__a31o_1 _06949_ (.A1(net548),
    .A2(net402),
    .A3(_00687_),
    .B1(_00686_),
    .X(_00813_));
 sky130_fd_sc_hd__nand4_1 _06950_ (.A(net548),
    .B(net447),
    .C(net394),
    .D(net378),
    .Y(_00814_));
 sky130_fd_sc_hd__a22o_1 _06951_ (.A1(net548),
    .A2(net394),
    .B1(net378),
    .B2(net447),
    .X(_00815_));
 sky130_fd_sc_hd__nand4_1 _06952_ (.A(net453),
    .B(net370),
    .C(_00814_),
    .D(_00815_),
    .Y(_00816_));
 sky130_fd_sc_hd__a22o_1 _06953_ (.A1(net453),
    .A2(net370),
    .B1(_00814_),
    .B2(_00815_),
    .X(_00817_));
 sky130_fd_sc_hd__nand3_1 _06954_ (.A(_00813_),
    .B(_00816_),
    .C(_00817_),
    .Y(_00818_));
 sky130_fd_sc_hd__a21o_1 _06955_ (.A1(_00816_),
    .A2(_00817_),
    .B1(_00813_),
    .X(_00819_));
 sky130_fd_sc_hd__nand3_1 _06956_ (.A(_00812_),
    .B(_00818_),
    .C(_00819_),
    .Y(_00820_));
 sky130_fd_sc_hd__a21o_1 _06957_ (.A1(_00818_),
    .A2(_00819_),
    .B1(_00812_),
    .X(_00821_));
 sky130_fd_sc_hd__a21bo_1 _06958_ (.A1(_00661_),
    .A2(_00670_),
    .B1_N(_00668_),
    .X(_00823_));
 sky130_fd_sc_hd__and3_1 _06959_ (.A(_00820_),
    .B(_00821_),
    .C(_00823_),
    .X(_00824_));
 sky130_fd_sc_hd__nand3_1 _06960_ (.A(_00820_),
    .B(_00821_),
    .C(_00823_),
    .Y(_00825_));
 sky130_fd_sc_hd__a21oi_1 _06961_ (.A1(_00820_),
    .A2(_00821_),
    .B1(_00823_),
    .Y(_00826_));
 sky130_fd_sc_hd__or3_2 _06962_ (.A(_00810_),
    .B(_00824_),
    .C(_00826_),
    .X(_00827_));
 sky130_fd_sc_hd__o21ai_1 _06963_ (.A1(_00824_),
    .A2(_00826_),
    .B1(_00810_),
    .Y(_00828_));
 sky130_fd_sc_hd__o211a_1 _06964_ (.A1(_00703_),
    .A2(_00705_),
    .B1(_00827_),
    .C1(_00828_),
    .X(_00829_));
 sky130_fd_sc_hd__a211oi_1 _06965_ (.A1(_00827_),
    .A2(_00828_),
    .B1(_00703_),
    .C1(_00705_),
    .Y(_00830_));
 sky130_fd_sc_hd__a211oi_1 _06966_ (.A1(_00675_),
    .A2(_00678_),
    .B1(_00829_),
    .C1(_00830_),
    .Y(_00831_));
 sky130_fd_sc_hd__o211a_1 _06967_ (.A1(_00829_),
    .A2(_00830_),
    .B1(_00675_),
    .C1(_00678_),
    .X(_00832_));
 sky130_fd_sc_hd__nand2_1 _06968_ (.A(net467),
    .B(net402),
    .Y(_00834_));
 sky130_fd_sc_hd__and4_1 _06969_ (.A(net387),
    .B(net416),
    .C(net303),
    .D(net408),
    .X(_00835_));
 sky130_fd_sc_hd__a22oi_1 _06970_ (.A1(net417),
    .A2(net301),
    .B1(net409),
    .B2(net387),
    .Y(_00836_));
 sky130_fd_sc_hd__nor2_1 _06971_ (.A(_00835_),
    .B(_00836_),
    .Y(_00837_));
 sky130_fd_sc_hd__xnor2_1 _06972_ (.A(_00834_),
    .B(_00837_),
    .Y(_00838_));
 sky130_fd_sc_hd__and4_1 _06973_ (.A(net185),
    .B(net429),
    .C(net181),
    .D(net172),
    .X(_00839_));
 sky130_fd_sc_hd__a22oi_1 _06974_ (.A1(net432),
    .A2(net181),
    .B1(net172),
    .B2(net185),
    .Y(_00840_));
 sky130_fd_sc_hd__and4bb_1 _06975_ (.A_N(_00839_),
    .B_N(_00840_),
    .C(net421),
    .D(net224),
    .X(_00841_));
 sky130_fd_sc_hd__o2bb2a_1 _06976_ (.A1_N(net425),
    .A2_N(net6),
    .B1(_00839_),
    .B2(_00840_),
    .X(_00842_));
 sky130_fd_sc_hd__nor2_1 _06977_ (.A(_00841_),
    .B(_00842_),
    .Y(_00843_));
 sky130_fd_sc_hd__nand2_1 _06978_ (.A(_00692_),
    .B(_00695_),
    .Y(_00845_));
 sky130_fd_sc_hd__and2_1 _06979_ (.A(_00843_),
    .B(_00845_),
    .X(_00846_));
 sky130_fd_sc_hd__xor2_1 _06980_ (.A(_00843_),
    .B(_00845_),
    .X(_00847_));
 sky130_fd_sc_hd__and2_1 _06981_ (.A(_00838_),
    .B(_00847_),
    .X(_00848_));
 sky130_fd_sc_hd__xnor2_1 _06982_ (.A(_00838_),
    .B(_00847_),
    .Y(_00849_));
 sky130_fd_sc_hd__a21oi_2 _06983_ (.A1(_00715_),
    .A2(_00717_),
    .B1(_00849_),
    .Y(_00850_));
 sky130_fd_sc_hd__inv_2 _06984_ (.A(_00850_),
    .Y(_00851_));
 sky130_fd_sc_hd__and3_1 _06985_ (.A(_00715_),
    .B(_00717_),
    .C(_00849_),
    .X(_00852_));
 sky130_fd_sc_hd__a211oi_1 _06986_ (.A1(_00698_),
    .A2(_00700_),
    .B1(_00850_),
    .C1(_00852_),
    .Y(_00853_));
 sky130_fd_sc_hd__a211o_1 _06987_ (.A1(_00698_),
    .A2(_00700_),
    .B1(_00850_),
    .C1(_00852_),
    .X(_00854_));
 sky130_fd_sc_hd__o211a_1 _06988_ (.A1(_00850_),
    .A2(_00852_),
    .B1(_00698_),
    .C1(_00700_),
    .X(_00855_));
 sky130_fd_sc_hd__o21ba_1 _06989_ (.A1(_00710_),
    .A2(_00712_),
    .B1_N(_00709_),
    .X(_00856_));
 sky130_fd_sc_hd__o21ba_1 _06990_ (.A1(_00720_),
    .A2(_00722_),
    .B1_N(_00719_),
    .X(_00857_));
 sky130_fd_sc_hd__nand2_1 _06991_ (.A(net195),
    .B(net164),
    .Y(_00858_));
 sky130_fd_sc_hd__and4_1 _06992_ (.A(net210),
    .B(net203),
    .C(net621),
    .D(net613),
    .X(_00859_));
 sky130_fd_sc_hd__a22oi_1 _06993_ (.A1(net203),
    .A2(net621),
    .B1(net613),
    .B2(net212),
    .Y(_00860_));
 sky130_fd_sc_hd__nor2_1 _06994_ (.A(_00859_),
    .B(_00860_),
    .Y(_00861_));
 sky130_fd_sc_hd__xnor2_1 _06995_ (.A(_00858_),
    .B(_00861_),
    .Y(_00862_));
 sky130_fd_sc_hd__nand2b_1 _06996_ (.A_N(_00857_),
    .B(_00862_),
    .Y(_00863_));
 sky130_fd_sc_hd__xnor2_1 _06997_ (.A(_00857_),
    .B(_00862_),
    .Y(_00864_));
 sky130_fd_sc_hd__nand2b_1 _06998_ (.A_N(_00856_),
    .B(_00864_),
    .Y(_00866_));
 sky130_fd_sc_hd__xnor2_1 _06999_ (.A(_00856_),
    .B(_00864_),
    .Y(_00867_));
 sky130_fd_sc_hd__nand2_1 _07000_ (.A(net218),
    .B(net597),
    .Y(_00868_));
 sky130_fd_sc_hd__and4_1 _07001_ (.A(net238),
    .B(net233),
    .C(net590),
    .D(net582),
    .X(_00869_));
 sky130_fd_sc_hd__a22oi_1 _07002_ (.A1(net233),
    .A2(net590),
    .B1(net582),
    .B2(net238),
    .Y(_00870_));
 sky130_fd_sc_hd__nor2_1 _07003_ (.A(_00869_),
    .B(_00870_),
    .Y(_00871_));
 sky130_fd_sc_hd__xnor2_1 _07004_ (.A(_00868_),
    .B(_00871_),
    .Y(_00872_));
 sky130_fd_sc_hd__and2_1 _07005_ (.A(net258),
    .B(net576),
    .X(_00873_));
 sky130_fd_sc_hd__nand4_1 _07006_ (.A(net437),
    .B(net345),
    .C(net568),
    .D(net562),
    .Y(_00874_));
 sky130_fd_sc_hd__a22o_1 _07007_ (.A1(net345),
    .A2(net568),
    .B1(net562),
    .B2(net437),
    .X(_00875_));
 sky130_fd_sc_hd__nand3_1 _07008_ (.A(_00873_),
    .B(_00874_),
    .C(_00875_),
    .Y(_00877_));
 sky130_fd_sc_hd__a21o_1 _07009_ (.A1(_00874_),
    .A2(_00875_),
    .B1(_00873_),
    .X(_00878_));
 sky130_fd_sc_hd__o21bai_1 _07010_ (.A1(_00725_),
    .A2(_00727_),
    .B1_N(_00726_),
    .Y(_00879_));
 sky130_fd_sc_hd__nand3_1 _07011_ (.A(_00877_),
    .B(_00878_),
    .C(_00879_),
    .Y(_00880_));
 sky130_fd_sc_hd__a21o_1 _07012_ (.A1(_00877_),
    .A2(_00878_),
    .B1(_00879_),
    .X(_00881_));
 sky130_fd_sc_hd__nand3_1 _07013_ (.A(_00872_),
    .B(_00880_),
    .C(_00881_),
    .Y(_00882_));
 sky130_fd_sc_hd__a21o_1 _07014_ (.A1(_00880_),
    .A2(_00881_),
    .B1(_00872_),
    .X(_00883_));
 sky130_fd_sc_hd__a21bo_1 _07015_ (.A1(_00723_),
    .A2(_00732_),
    .B1_N(_00731_),
    .X(_00884_));
 sky130_fd_sc_hd__nand3_2 _07016_ (.A(_00882_),
    .B(_00883_),
    .C(_00884_),
    .Y(_00885_));
 sky130_fd_sc_hd__a21o_1 _07017_ (.A1(_00882_),
    .A2(_00883_),
    .B1(_00884_),
    .X(_00886_));
 sky130_fd_sc_hd__and3_1 _07018_ (.A(_00867_),
    .B(_00885_),
    .C(_00886_),
    .X(_00888_));
 sky130_fd_sc_hd__nand3_1 _07019_ (.A(_00867_),
    .B(_00885_),
    .C(_00886_),
    .Y(_00889_));
 sky130_fd_sc_hd__a21oi_1 _07020_ (.A1(_00885_),
    .A2(_00886_),
    .B1(_00867_),
    .Y(_00890_));
 sky130_fd_sc_hd__a211oi_2 _07021_ (.A1(_00737_),
    .A2(_00740_),
    .B1(_00888_),
    .C1(_00890_),
    .Y(_00891_));
 sky130_fd_sc_hd__o211a_1 _07022_ (.A1(_00888_),
    .A2(_00890_),
    .B1(_00737_),
    .C1(_00740_),
    .X(_00892_));
 sky130_fd_sc_hd__nor4_1 _07023_ (.A(_00853_),
    .B(_00855_),
    .C(_00891_),
    .D(_00892_),
    .Y(_00893_));
 sky130_fd_sc_hd__o22a_1 _07024_ (.A1(_00853_),
    .A2(_00855_),
    .B1(_00891_),
    .B2(_00892_),
    .X(_00894_));
 sky130_fd_sc_hd__a211o_1 _07025_ (.A1(_00742_),
    .A2(_00744_),
    .B1(net146),
    .C1(_00894_),
    .X(_00895_));
 sky130_fd_sc_hd__o211ai_1 _07026_ (.A1(net146),
    .A2(_00894_),
    .B1(_00742_),
    .C1(_00744_),
    .Y(_00896_));
 sky130_fd_sc_hd__or4bb_2 _07027_ (.A(_00831_),
    .B(_00832_),
    .C_N(_00895_),
    .D_N(_00896_),
    .X(_00897_));
 sky130_fd_sc_hd__a2bb2o_1 _07028_ (.A1_N(_00831_),
    .A2_N(_00832_),
    .B1(_00895_),
    .B2(_00896_),
    .X(_00899_));
 sky130_fd_sc_hd__o211a_2 _07029_ (.A1(_00747_),
    .A2(_00749_),
    .B1(_00897_),
    .C1(_00899_),
    .X(_00900_));
 sky130_fd_sc_hd__a211oi_1 _07030_ (.A1(_00897_),
    .A2(_00899_),
    .B1(_00747_),
    .C1(_00749_),
    .Y(_00901_));
 sky130_fd_sc_hd__nor3_1 _07031_ (.A(_00794_),
    .B(_00900_),
    .C(_00901_),
    .Y(_00902_));
 sky130_fd_sc_hd__or3_1 _07032_ (.A(_00794_),
    .B(_00900_),
    .C(_00901_),
    .X(_00903_));
 sky130_fd_sc_hd__o21ai_1 _07033_ (.A1(_00900_),
    .A2(_00901_),
    .B1(_00794_),
    .Y(_00904_));
 sky130_fd_sc_hd__o211a_1 _07034_ (.A1(_00751_),
    .A2(_00753_),
    .B1(_00903_),
    .C1(_00904_),
    .X(_00905_));
 sky130_fd_sc_hd__a211oi_1 _07035_ (.A1(_00903_),
    .A2(_00904_),
    .B1(_00751_),
    .C1(_00753_),
    .Y(_00906_));
 sky130_fd_sc_hd__nor3_1 _07036_ (.A(_00641_),
    .B(_00905_),
    .C(_00906_),
    .Y(_00907_));
 sky130_fd_sc_hd__o21a_1 _07037_ (.A1(_00905_),
    .A2(_00906_),
    .B1(_00641_),
    .X(_00908_));
 sky130_fd_sc_hd__a211o_1 _07038_ (.A1(_00756_),
    .A2(_00759_),
    .B1(net130),
    .C1(_00908_),
    .X(_00910_));
 sky130_fd_sc_hd__o211ai_1 _07039_ (.A1(net130),
    .A2(_00908_),
    .B1(_00756_),
    .C1(_00759_),
    .Y(_00911_));
 sky130_fd_sc_hd__a21oi_1 _07040_ (.A1(_00910_),
    .A2(_00911_),
    .B1(_00761_),
    .Y(_00912_));
 sky130_fd_sc_hd__inv_2 _07041_ (.A(_00912_),
    .Y(_00913_));
 sky130_fd_sc_hd__and3_1 _07042_ (.A(_00761_),
    .B(_00910_),
    .C(_00911_),
    .X(_00914_));
 sky130_fd_sc_hd__nor2_1 _07043_ (.A(_00912_),
    .B(_00914_),
    .Y(_00915_));
 sky130_fd_sc_hd__o21ba_1 _07044_ (.A1(_00765_),
    .A2(_00773_),
    .B1_N(_00764_),
    .X(_00916_));
 sky130_fd_sc_hd__xnor2_1 _07045_ (.A(_00915_),
    .B(_00916_),
    .Y(net82));
 sky130_fd_sc_hd__or2_1 _07046_ (.A(_00829_),
    .B(_00831_),
    .X(_00917_));
 sky130_fd_sc_hd__a21oi_1 _07047_ (.A1(_00799_),
    .A2(_00808_),
    .B1(_00807_),
    .Y(_00918_));
 sky130_fd_sc_hd__a31o_1 _07048_ (.A1(net518),
    .A2(net318),
    .A3(_00797_),
    .B1(_00796_),
    .X(_00920_));
 sky130_fd_sc_hd__nand4_1 _07049_ (.A(net518),
    .B(net602),
    .C(net310),
    .D(net296),
    .Y(_00921_));
 sky130_fd_sc_hd__a22o_1 _07050_ (.A1(net518),
    .A2(net311),
    .B1(net296),
    .B2(net602),
    .X(_00922_));
 sky130_fd_sc_hd__nand2_1 _07051_ (.A(net628),
    .B(net288),
    .Y(_00923_));
 sky130_fd_sc_hd__nand3b_1 _07052_ (.A_N(_00923_),
    .B(_00922_),
    .C(_00921_),
    .Y(_00924_));
 sky130_fd_sc_hd__a21bo_1 _07053_ (.A1(_00921_),
    .A2(_00922_),
    .B1_N(_00923_),
    .X(_00925_));
 sky130_fd_sc_hd__and3_1 _07054_ (.A(_00920_),
    .B(_00924_),
    .C(_00925_),
    .X(_00926_));
 sky130_fd_sc_hd__a21o_1 _07055_ (.A1(_00924_),
    .A2(_00925_),
    .B1(_00920_),
    .X(_00927_));
 sky130_fd_sc_hd__and2b_1 _07056_ (.A_N(_00926_),
    .B(_00927_),
    .X(_00928_));
 sky130_fd_sc_hd__xnor2_1 _07057_ (.A(_00777_),
    .B(_00928_),
    .Y(_00929_));
 sky130_fd_sc_hd__nor2_1 _07058_ (.A(_00918_),
    .B(_00929_),
    .Y(_00931_));
 sky130_fd_sc_hd__xor2_1 _07059_ (.A(_00918_),
    .B(_00929_),
    .X(_00932_));
 sky130_fd_sc_hd__xnor2_1 _07060_ (.A(_00780_),
    .B(_00932_),
    .Y(_00933_));
 sky130_fd_sc_hd__a21o_1 _07061_ (.A1(_00783_),
    .A2(_00785_),
    .B1(_00933_),
    .X(_00934_));
 sky130_fd_sc_hd__nand3_1 _07062_ (.A(_00783_),
    .B(_00785_),
    .C(_00933_),
    .Y(_00935_));
 sky130_fd_sc_hd__nand2_1 _07063_ (.A(_00934_),
    .B(_00935_),
    .Y(_00936_));
 sky130_fd_sc_hd__nand2b_1 _07064_ (.A_N(_00936_),
    .B(_00917_),
    .Y(_00937_));
 sky130_fd_sc_hd__xnor2_1 _07065_ (.A(_00917_),
    .B(_00936_),
    .Y(_00938_));
 sky130_fd_sc_hd__nand2_1 _07066_ (.A(_00787_),
    .B(_00938_),
    .Y(_00939_));
 sky130_fd_sc_hd__xnor2_1 _07067_ (.A(_00787_),
    .B(_00938_),
    .Y(_00940_));
 sky130_fd_sc_hd__nand2_1 _07068_ (.A(net498),
    .B(net318),
    .Y(_00941_));
 sky130_fd_sc_hd__and4_1 _07069_ (.A(net484),
    .B(net490),
    .C(net332),
    .D(net325),
    .X(_00942_));
 sky130_fd_sc_hd__a22oi_1 _07070_ (.A1(net484),
    .A2(net332),
    .B1(net325),
    .B2(net490),
    .Y(_00943_));
 sky130_fd_sc_hd__nor2_1 _07071_ (.A(_00942_),
    .B(_00943_),
    .Y(_00944_));
 sky130_fd_sc_hd__xnor2_1 _07072_ (.A(_00941_),
    .B(_00944_),
    .Y(_00945_));
 sky130_fd_sc_hd__and4_1 _07073_ (.A(net461),
    .B(net454),
    .C(net363),
    .D(net355),
    .X(_00946_));
 sky130_fd_sc_hd__a22oi_1 _07074_ (.A1(net454),
    .A2(net363),
    .B1(net355),
    .B2(net461),
    .Y(_00947_));
 sky130_fd_sc_hd__and4bb_1 _07075_ (.A_N(_00946_),
    .B_N(_00947_),
    .C(net476),
    .D(net340),
    .X(_00948_));
 sky130_fd_sc_hd__o2bb2a_1 _07076_ (.A1_N(net476),
    .A2_N(net340),
    .B1(_00946_),
    .B2(_00947_),
    .X(_00949_));
 sky130_fd_sc_hd__o21ba_1 _07077_ (.A1(_00801_),
    .A2(_00803_),
    .B1_N(_00802_),
    .X(_00950_));
 sky130_fd_sc_hd__nor3_1 _07078_ (.A(_00948_),
    .B(_00949_),
    .C(_00950_),
    .Y(_00952_));
 sky130_fd_sc_hd__o21a_1 _07079_ (.A1(_00948_),
    .A2(_00949_),
    .B1(_00950_),
    .X(_00953_));
 sky130_fd_sc_hd__nor2_1 _07080_ (.A(_00952_),
    .B(_00953_),
    .Y(_00954_));
 sky130_fd_sc_hd__xnor2_1 _07081_ (.A(_00945_),
    .B(_00954_),
    .Y(_00955_));
 sky130_fd_sc_hd__nand2_1 _07082_ (.A(_00814_),
    .B(_00816_),
    .Y(_00956_));
 sky130_fd_sc_hd__o21ba_1 _07083_ (.A1(_00834_),
    .A2(_00836_),
    .B1_N(_00835_),
    .X(_00957_));
 sky130_fd_sc_hd__nand2_1 _07084_ (.A(net448),
    .B(net370),
    .Y(_00958_));
 sky130_fd_sc_hd__and4_1 _07085_ (.A(net549),
    .B(net468),
    .C(net392),
    .D(net376),
    .X(_00959_));
 sky130_fd_sc_hd__a22oi_1 _07086_ (.A1(net468),
    .A2(net394),
    .B1(net376),
    .B2(net549),
    .Y(_00960_));
 sky130_fd_sc_hd__nor2_1 _07087_ (.A(_00959_),
    .B(_00960_),
    .Y(_00961_));
 sky130_fd_sc_hd__xnor2_1 _07088_ (.A(_00958_),
    .B(_00961_),
    .Y(_00963_));
 sky130_fd_sc_hd__nand2b_1 _07089_ (.A_N(_00957_),
    .B(_00963_),
    .Y(_00964_));
 sky130_fd_sc_hd__xnor2_1 _07090_ (.A(_00957_),
    .B(_00963_),
    .Y(_00965_));
 sky130_fd_sc_hd__nand2_1 _07091_ (.A(_00956_),
    .B(_00965_),
    .Y(_00966_));
 sky130_fd_sc_hd__xnor2_1 _07092_ (.A(_00956_),
    .B(_00965_),
    .Y(_00967_));
 sky130_fd_sc_hd__a21oi_1 _07093_ (.A1(_00818_),
    .A2(_00820_),
    .B1(_00967_),
    .Y(_00968_));
 sky130_fd_sc_hd__inv_2 _07094_ (.A(_00968_),
    .Y(_00969_));
 sky130_fd_sc_hd__and3_1 _07095_ (.A(_00818_),
    .B(_00820_),
    .C(_00967_),
    .X(_00970_));
 sky130_fd_sc_hd__nor3_1 _07096_ (.A(_00955_),
    .B(_00968_),
    .C(_00970_),
    .Y(_00971_));
 sky130_fd_sc_hd__inv_2 _07097_ (.A(_00971_),
    .Y(_00972_));
 sky130_fd_sc_hd__o21a_1 _07098_ (.A1(_00968_),
    .A2(_00970_),
    .B1(_00955_),
    .X(_00974_));
 sky130_fd_sc_hd__a211oi_2 _07099_ (.A1(_00851_),
    .A2(_00854_),
    .B1(net153),
    .C1(_00974_),
    .Y(_00975_));
 sky130_fd_sc_hd__o211a_1 _07100_ (.A1(net153),
    .A2(_00974_),
    .B1(_00851_),
    .C1(_00854_),
    .X(_00976_));
 sky130_fd_sc_hd__a211oi_2 _07101_ (.A1(_00825_),
    .A2(_00827_),
    .B1(_00975_),
    .C1(_00976_),
    .Y(_00977_));
 sky130_fd_sc_hd__o211a_1 _07102_ (.A1(_00975_),
    .A2(_00976_),
    .B1(_00825_),
    .C1(_00827_),
    .X(_00978_));
 sky130_fd_sc_hd__nand2_1 _07103_ (.A(net386),
    .B(net401),
    .Y(_00979_));
 sky130_fd_sc_hd__and4_1 _07104_ (.A(net416),
    .B(net301),
    .C(net408),
    .D(net225),
    .X(_00980_));
 sky130_fd_sc_hd__a22oi_1 _07105_ (.A1(net301),
    .A2(net408),
    .B1(net225),
    .B2(net416),
    .Y(_00981_));
 sky130_fd_sc_hd__nor2_1 _07106_ (.A(_00980_),
    .B(_00981_),
    .Y(_00982_));
 sky130_fd_sc_hd__xnor2_1 _07107_ (.A(_00979_),
    .B(_00982_),
    .Y(_00983_));
 sky130_fd_sc_hd__nand2_1 _07108_ (.A(net425),
    .B(net180),
    .Y(_00985_));
 sky130_fd_sc_hd__and4_1 _07109_ (.A(net185),
    .B(net429),
    .C(net173),
    .D(net165),
    .X(_00986_));
 sky130_fd_sc_hd__a22oi_1 _07110_ (.A1(net429),
    .A2(net172),
    .B1(net164),
    .B2(net185),
    .Y(_00987_));
 sky130_fd_sc_hd__nor2_1 _07111_ (.A(_00986_),
    .B(_00987_),
    .Y(_00988_));
 sky130_fd_sc_hd__xnor2_1 _07112_ (.A(_00985_),
    .B(_00988_),
    .Y(_00989_));
 sky130_fd_sc_hd__nor2_1 _07113_ (.A(_00839_),
    .B(_00841_),
    .Y(_00990_));
 sky130_fd_sc_hd__and2b_1 _07114_ (.A_N(_00990_),
    .B(_00989_),
    .X(_00991_));
 sky130_fd_sc_hd__xnor2_1 _07115_ (.A(_00989_),
    .B(_00990_),
    .Y(_00992_));
 sky130_fd_sc_hd__and2_1 _07116_ (.A(_00983_),
    .B(_00992_),
    .X(_00993_));
 sky130_fd_sc_hd__xnor2_1 _07117_ (.A(_00983_),
    .B(_00992_),
    .Y(_00994_));
 sky130_fd_sc_hd__a21oi_1 _07118_ (.A1(_00863_),
    .A2(_00866_),
    .B1(_00994_),
    .Y(_00996_));
 sky130_fd_sc_hd__a21o_1 _07119_ (.A1(_00863_),
    .A2(_00866_),
    .B1(_00994_),
    .X(_00997_));
 sky130_fd_sc_hd__nand3_1 _07120_ (.A(_00863_),
    .B(_00866_),
    .C(_00994_),
    .Y(_00998_));
 sky130_fd_sc_hd__o211a_1 _07121_ (.A1(_00846_),
    .A2(_00848_),
    .B1(_00997_),
    .C1(_00998_),
    .X(_00999_));
 sky130_fd_sc_hd__a211oi_1 _07122_ (.A1(_00997_),
    .A2(_00998_),
    .B1(_00846_),
    .C1(_00848_),
    .Y(_01000_));
 sky130_fd_sc_hd__o21ba_1 _07123_ (.A1(_00858_),
    .A2(_00860_),
    .B1_N(_00859_),
    .X(_01001_));
 sky130_fd_sc_hd__o21ba_1 _07124_ (.A1(_00868_),
    .A2(_00870_),
    .B1_N(_00869_),
    .X(_01002_));
 sky130_fd_sc_hd__nand2_1 _07125_ (.A(net193),
    .B(net620),
    .Y(_01003_));
 sky130_fd_sc_hd__and4_1 _07126_ (.A(net210),
    .B(net201),
    .C(net612),
    .D(net596),
    .X(_01004_));
 sky130_fd_sc_hd__a22oi_1 _07127_ (.A1(net201),
    .A2(net612),
    .B1(net596),
    .B2(net210),
    .Y(_01005_));
 sky130_fd_sc_hd__nor2_1 _07128_ (.A(_01004_),
    .B(_01005_),
    .Y(_01007_));
 sky130_fd_sc_hd__xnor2_1 _07129_ (.A(_01003_),
    .B(_01007_),
    .Y(_01008_));
 sky130_fd_sc_hd__nand2b_1 _07130_ (.A_N(_01002_),
    .B(_01008_),
    .Y(_01009_));
 sky130_fd_sc_hd__xnor2_1 _07131_ (.A(_01002_),
    .B(_01008_),
    .Y(_01010_));
 sky130_fd_sc_hd__nand2b_1 _07132_ (.A_N(_01001_),
    .B(_01010_),
    .Y(_01011_));
 sky130_fd_sc_hd__xnor2_1 _07133_ (.A(_01001_),
    .B(_01010_),
    .Y(_01012_));
 sky130_fd_sc_hd__nand2_1 _07134_ (.A(net218),
    .B(net589),
    .Y(_01013_));
 sky130_fd_sc_hd__and4_1 _07135_ (.A(net238),
    .B(net229),
    .C(net581),
    .D(net575),
    .X(_01014_));
 sky130_fd_sc_hd__a22oi_1 _07136_ (.A1(net229),
    .A2(net582),
    .B1(net576),
    .B2(net238),
    .Y(_01015_));
 sky130_fd_sc_hd__nor2_1 _07137_ (.A(_01014_),
    .B(_01015_),
    .Y(_01016_));
 sky130_fd_sc_hd__xnor2_1 _07138_ (.A(_01013_),
    .B(_01016_),
    .Y(_01018_));
 sky130_fd_sc_hd__nand2_1 _07139_ (.A(net257),
    .B(net568),
    .Y(_01019_));
 sky130_fd_sc_hd__and4_1 _07140_ (.A(net436),
    .B(net343),
    .C(net562),
    .D(net554),
    .X(_01020_));
 sky130_fd_sc_hd__a22oi_2 _07141_ (.A1(net346),
    .A2(net562),
    .B1(net554),
    .B2(net436),
    .Y(_01021_));
 sky130_fd_sc_hd__or3_1 _07142_ (.A(_01019_),
    .B(_01020_),
    .C(_01021_),
    .X(_01022_));
 sky130_fd_sc_hd__o21ai_1 _07143_ (.A1(_01020_),
    .A2(_01021_),
    .B1(_01019_),
    .Y(_01023_));
 sky130_fd_sc_hd__a21bo_1 _07144_ (.A1(_00873_),
    .A2(_00875_),
    .B1_N(_00874_),
    .X(_01024_));
 sky130_fd_sc_hd__nand3_1 _07145_ (.A(_01022_),
    .B(_01023_),
    .C(_01024_),
    .Y(_01025_));
 sky130_fd_sc_hd__a21o_1 _07146_ (.A1(_01022_),
    .A2(_01023_),
    .B1(_01024_),
    .X(_01026_));
 sky130_fd_sc_hd__nand3_1 _07147_ (.A(_01018_),
    .B(_01025_),
    .C(_01026_),
    .Y(_01027_));
 sky130_fd_sc_hd__a21o_1 _07148_ (.A1(_01025_),
    .A2(_01026_),
    .B1(_01018_),
    .X(_01029_));
 sky130_fd_sc_hd__a21bo_1 _07149_ (.A1(_00872_),
    .A2(_00881_),
    .B1_N(_00880_),
    .X(_01030_));
 sky130_fd_sc_hd__nand3_2 _07150_ (.A(_01027_),
    .B(_01029_),
    .C(_01030_),
    .Y(_01031_));
 sky130_fd_sc_hd__a21o_1 _07151_ (.A1(_01027_),
    .A2(_01029_),
    .B1(_01030_),
    .X(_01032_));
 sky130_fd_sc_hd__and3_1 _07152_ (.A(_01012_),
    .B(_01031_),
    .C(_01032_),
    .X(_01033_));
 sky130_fd_sc_hd__nand3_1 _07153_ (.A(_01012_),
    .B(_01031_),
    .C(_01032_),
    .Y(_01034_));
 sky130_fd_sc_hd__a21oi_1 _07154_ (.A1(_01031_),
    .A2(_01032_),
    .B1(_01012_),
    .Y(_01035_));
 sky130_fd_sc_hd__a211o_1 _07155_ (.A1(_00885_),
    .A2(_00889_),
    .B1(_01033_),
    .C1(_01035_),
    .X(_01036_));
 sky130_fd_sc_hd__o211ai_1 _07156_ (.A1(_01033_),
    .A2(_01035_),
    .B1(_00885_),
    .C1(_00889_),
    .Y(_01037_));
 sky130_fd_sc_hd__or4bb_2 _07157_ (.A(_00999_),
    .B(_01000_),
    .C_N(_01036_),
    .D_N(_01037_),
    .X(_01038_));
 sky130_fd_sc_hd__a2bb2o_1 _07158_ (.A1_N(_00999_),
    .A2_N(_01000_),
    .B1(_01036_),
    .B2(_01037_),
    .X(_01040_));
 sky130_fd_sc_hd__o211a_2 _07159_ (.A1(_00891_),
    .A2(_00893_),
    .B1(_01038_),
    .C1(_01040_),
    .X(_01041_));
 sky130_fd_sc_hd__a211oi_1 _07160_ (.A1(_01038_),
    .A2(_01040_),
    .B1(_00891_),
    .C1(_00893_),
    .Y(_01042_));
 sky130_fd_sc_hd__nor4_1 _07161_ (.A(_00977_),
    .B(_00978_),
    .C(_01041_),
    .D(_01042_),
    .Y(_01043_));
 sky130_fd_sc_hd__o22a_1 _07162_ (.A1(_00977_),
    .A2(_00978_),
    .B1(_01041_),
    .B2(_01042_),
    .X(_01044_));
 sky130_fd_sc_hd__a211oi_2 _07163_ (.A1(_00895_),
    .A2(_00897_),
    .B1(net140),
    .C1(_01044_),
    .Y(_01045_));
 sky130_fd_sc_hd__o211a_1 _07164_ (.A1(net140),
    .A2(_01044_),
    .B1(_00895_),
    .C1(_00897_),
    .X(_01046_));
 sky130_fd_sc_hd__nor3_1 _07165_ (.A(_00940_),
    .B(_01045_),
    .C(_01046_),
    .Y(_01047_));
 sky130_fd_sc_hd__or3_2 _07166_ (.A(_00940_),
    .B(_01045_),
    .C(_01046_),
    .X(_01048_));
 sky130_fd_sc_hd__o21ai_2 _07167_ (.A1(_01045_),
    .A2(_01046_),
    .B1(_00940_),
    .Y(_01049_));
 sky130_fd_sc_hd__o211ai_4 _07168_ (.A1(_00900_),
    .A2(net133),
    .B1(_01048_),
    .C1(_01049_),
    .Y(_01051_));
 sky130_fd_sc_hd__a211o_1 _07169_ (.A1(_01048_),
    .A2(_01049_),
    .B1(_00900_),
    .C1(_00902_),
    .X(_01052_));
 sky130_fd_sc_hd__o211ai_4 _07170_ (.A1(_00791_),
    .A2(_00793_),
    .B1(_01051_),
    .C1(_01052_),
    .Y(_01053_));
 sky130_fd_sc_hd__a211o_1 _07171_ (.A1(_01051_),
    .A2(_01052_),
    .B1(_00791_),
    .C1(_00793_),
    .X(_01054_));
 sky130_fd_sc_hd__o211a_1 _07172_ (.A1(_00905_),
    .A2(_00907_),
    .B1(_01053_),
    .C1(_01054_),
    .X(_01055_));
 sky130_fd_sc_hd__a211oi_1 _07173_ (.A1(_01053_),
    .A2(_01054_),
    .B1(_00905_),
    .C1(_00907_),
    .Y(_01056_));
 sky130_fd_sc_hd__or2_1 _07174_ (.A(_01055_),
    .B(_01056_),
    .X(_01057_));
 sky130_fd_sc_hd__nor2_1 _07175_ (.A(_00910_),
    .B(_01057_),
    .Y(_01058_));
 sky130_fd_sc_hd__xnor2_1 _07176_ (.A(_00910_),
    .B(_01057_),
    .Y(_01059_));
 sky130_fd_sc_hd__a21oi_1 _07177_ (.A1(_00764_),
    .A2(_00913_),
    .B1(_00914_),
    .Y(_01060_));
 sky130_fd_sc_hd__or3_1 _07178_ (.A(_00765_),
    .B(_00912_),
    .C(_00914_),
    .X(_01062_));
 sky130_fd_sc_hd__o21a_1 _07179_ (.A1(_00773_),
    .A2(_01062_),
    .B1(_01060_),
    .X(_01063_));
 sky130_fd_sc_hd__nor2_1 _07180_ (.A(_01059_),
    .B(_01063_),
    .Y(_01064_));
 sky130_fd_sc_hd__xor2_1 _07181_ (.A(_01059_),
    .B(_01063_),
    .X(net83));
 sky130_fd_sc_hd__a21o_1 _07182_ (.A1(_00777_),
    .A2(_00927_),
    .B1(_00926_),
    .X(_01065_));
 sky130_fd_sc_hd__a21oi_1 _07183_ (.A1(_00945_),
    .A2(_00954_),
    .B1(_00952_),
    .Y(_01066_));
 sky130_fd_sc_hd__nand2_1 _07184_ (.A(_00921_),
    .B(_00924_),
    .Y(_01067_));
 sky130_fd_sc_hd__o21ba_1 _07185_ (.A1(_00941_),
    .A2(_00943_),
    .B1_N(_00942_),
    .X(_01068_));
 sky130_fd_sc_hd__and4_1 _07186_ (.A(net496),
    .B(net517),
    .C(net310),
    .D(net296),
    .X(_01069_));
 sky130_fd_sc_hd__a22oi_1 _07187_ (.A1(net498),
    .A2(net310),
    .B1(net296),
    .B2(net517),
    .Y(_01070_));
 sky130_fd_sc_hd__o2bb2a_1 _07188_ (.A1_N(net603),
    .A2_N(net288),
    .B1(_01069_),
    .B2(_01070_),
    .X(_01072_));
 sky130_fd_sc_hd__and4bb_1 _07189_ (.A_N(_01069_),
    .B_N(_01070_),
    .C(net603),
    .D(net288),
    .X(_01073_));
 sky130_fd_sc_hd__nor2_1 _07190_ (.A(_01072_),
    .B(_01073_),
    .Y(_01074_));
 sky130_fd_sc_hd__or3_1 _07191_ (.A(_01068_),
    .B(_01072_),
    .C(_01073_),
    .X(_01075_));
 sky130_fd_sc_hd__xnor2_1 _07192_ (.A(_01068_),
    .B(_01074_),
    .Y(_01076_));
 sky130_fd_sc_hd__nand2_1 _07193_ (.A(_01067_),
    .B(_01076_),
    .Y(_01077_));
 sky130_fd_sc_hd__xor2_1 _07194_ (.A(_01067_),
    .B(_01076_),
    .X(_01078_));
 sky130_fd_sc_hd__and2b_1 _07195_ (.A_N(_01066_),
    .B(_01078_),
    .X(_01079_));
 sky130_fd_sc_hd__xnor2_1 _07196_ (.A(_01066_),
    .B(_01078_),
    .Y(_01080_));
 sky130_fd_sc_hd__and2_1 _07197_ (.A(_01065_),
    .B(_01080_),
    .X(_01081_));
 sky130_fd_sc_hd__xnor2_1 _07198_ (.A(_01065_),
    .B(_01080_),
    .Y(_01083_));
 sky130_fd_sc_hd__a21oi_1 _07199_ (.A1(_00780_),
    .A2(_00932_),
    .B1(_00931_),
    .Y(_01084_));
 sky130_fd_sc_hd__or2_1 _07200_ (.A(_01083_),
    .B(_01084_),
    .X(_01085_));
 sky130_fd_sc_hd__xnor2_1 _07201_ (.A(_01083_),
    .B(_01084_),
    .Y(_01086_));
 sky130_fd_sc_hd__nand2_1 _07202_ (.A(net628),
    .B(net282),
    .Y(_01087_));
 sky130_fd_sc_hd__or2_1 _07203_ (.A(_01086_),
    .B(_01087_),
    .X(_01088_));
 sky130_fd_sc_hd__xor2_1 _07204_ (.A(_01086_),
    .B(_01087_),
    .X(_01089_));
 sky130_fd_sc_hd__nor3_1 _07205_ (.A(_00975_),
    .B(_00977_),
    .C(_01089_),
    .Y(_01090_));
 sky130_fd_sc_hd__o21a_1 _07206_ (.A1(_00975_),
    .A2(_00977_),
    .B1(_01089_),
    .X(_01091_));
 sky130_fd_sc_hd__o21ai_1 _07207_ (.A1(_01090_),
    .A2(_01091_),
    .B1(_00934_),
    .Y(_01092_));
 sky130_fd_sc_hd__or3_1 _07208_ (.A(_00934_),
    .B(_01090_),
    .C(_01091_),
    .X(_01094_));
 sky130_fd_sc_hd__and4_1 _07209_ (.A(net484),
    .B(net476),
    .C(net332),
    .D(net325),
    .X(_01095_));
 sky130_fd_sc_hd__a22oi_1 _07210_ (.A1(net476),
    .A2(net332),
    .B1(net325),
    .B2(net484),
    .Y(_01096_));
 sky130_fd_sc_hd__and4bb_1 _07211_ (.A_N(_01095_),
    .B_N(_01096_),
    .C(net490),
    .D(net318),
    .X(_01097_));
 sky130_fd_sc_hd__o2bb2a_1 _07212_ (.A1_N(net490),
    .A2_N(net48),
    .B1(_01095_),
    .B2(_01096_),
    .X(_01098_));
 sky130_fd_sc_hd__nor2_1 _07213_ (.A(_01097_),
    .B(_01098_),
    .Y(_01099_));
 sky130_fd_sc_hd__nand2_1 _07214_ (.A(net461),
    .B(net339),
    .Y(_01100_));
 sky130_fd_sc_hd__and4_1 _07215_ (.A(net455),
    .B(net448),
    .C(net361),
    .D(net353),
    .X(_01101_));
 sky130_fd_sc_hd__a22oi_1 _07216_ (.A1(net448),
    .A2(net361),
    .B1(net353),
    .B2(net455),
    .Y(_01102_));
 sky130_fd_sc_hd__nor2_1 _07217_ (.A(_01101_),
    .B(_01102_),
    .Y(_01103_));
 sky130_fd_sc_hd__xnor2_1 _07218_ (.A(_01100_),
    .B(_01103_),
    .Y(_01105_));
 sky130_fd_sc_hd__nor2_1 _07219_ (.A(_00946_),
    .B(_00948_),
    .Y(_01106_));
 sky130_fd_sc_hd__and2b_1 _07220_ (.A_N(_01106_),
    .B(_01105_),
    .X(_01107_));
 sky130_fd_sc_hd__xnor2_1 _07221_ (.A(_01105_),
    .B(_01106_),
    .Y(_01108_));
 sky130_fd_sc_hd__and2_1 _07222_ (.A(_01099_),
    .B(_01108_),
    .X(_01109_));
 sky130_fd_sc_hd__nor2_1 _07223_ (.A(_01099_),
    .B(_01108_),
    .Y(_01110_));
 sky130_fd_sc_hd__or2_1 _07224_ (.A(_01109_),
    .B(_01110_),
    .X(_01111_));
 sky130_fd_sc_hd__a31o_1 _07225_ (.A1(net448),
    .A2(net369),
    .A3(_00961_),
    .B1(_00959_),
    .X(_01112_));
 sky130_fd_sc_hd__o21ba_1 _07226_ (.A1(_00979_),
    .A2(_00981_),
    .B1_N(_00980_),
    .X(_01113_));
 sky130_fd_sc_hd__nand2_1 _07227_ (.A(net549),
    .B(net369),
    .Y(_01114_));
 sky130_fd_sc_hd__and4_1 _07228_ (.A(net468),
    .B(net386),
    .C(net392),
    .D(net376),
    .X(_01116_));
 sky130_fd_sc_hd__a22oi_1 _07229_ (.A1(net386),
    .A2(net392),
    .B1(net376),
    .B2(net468),
    .Y(_01117_));
 sky130_fd_sc_hd__nor2_1 _07230_ (.A(_01116_),
    .B(_01117_),
    .Y(_01118_));
 sky130_fd_sc_hd__xnor2_1 _07231_ (.A(_01114_),
    .B(_01118_),
    .Y(_01119_));
 sky130_fd_sc_hd__nand2b_1 _07232_ (.A_N(_01113_),
    .B(_01119_),
    .Y(_01120_));
 sky130_fd_sc_hd__xnor2_1 _07233_ (.A(_01113_),
    .B(_01119_),
    .Y(_01121_));
 sky130_fd_sc_hd__nand2_1 _07234_ (.A(_01112_),
    .B(_01121_),
    .Y(_01122_));
 sky130_fd_sc_hd__xnor2_1 _07235_ (.A(_01112_),
    .B(_01121_),
    .Y(_01123_));
 sky130_fd_sc_hd__a21o_1 _07236_ (.A1(_00964_),
    .A2(_00966_),
    .B1(_01123_),
    .X(_01124_));
 sky130_fd_sc_hd__nand3_1 _07237_ (.A(_00964_),
    .B(_00966_),
    .C(_01123_),
    .Y(_01125_));
 sky130_fd_sc_hd__nand3b_2 _07238_ (.A_N(_01111_),
    .B(_01124_),
    .C(_01125_),
    .Y(_01127_));
 sky130_fd_sc_hd__a21bo_1 _07239_ (.A1(_01124_),
    .A2(_01125_),
    .B1_N(_01111_),
    .X(_01128_));
 sky130_fd_sc_hd__o211a_1 _07240_ (.A1(_00996_),
    .A2(_00999_),
    .B1(_01127_),
    .C1(_01128_),
    .X(_01129_));
 sky130_fd_sc_hd__a211oi_1 _07241_ (.A1(_01127_),
    .A2(_01128_),
    .B1(_00996_),
    .C1(_00999_),
    .Y(_01130_));
 sky130_fd_sc_hd__a211oi_2 _07242_ (.A1(_00969_),
    .A2(_00972_),
    .B1(_01129_),
    .C1(_01130_),
    .Y(_01131_));
 sky130_fd_sc_hd__o211a_1 _07243_ (.A1(_01129_),
    .A2(_01130_),
    .B1(_00969_),
    .C1(_00972_),
    .X(_01132_));
 sky130_fd_sc_hd__nand2_1 _07244_ (.A(net301),
    .B(net401),
    .Y(_01133_));
 sky130_fd_sc_hd__and4_1 _07245_ (.A(net416),
    .B(net408),
    .C(net225),
    .D(net180),
    .X(_01134_));
 sky130_fd_sc_hd__a22oi_1 _07246_ (.A1(net408),
    .A2(net225),
    .B1(net180),
    .B2(net416),
    .Y(_01135_));
 sky130_fd_sc_hd__nor2_1 _07247_ (.A(_01134_),
    .B(_01135_),
    .Y(_01136_));
 sky130_fd_sc_hd__xnor2_1 _07248_ (.A(_01133_),
    .B(_01136_),
    .Y(_01138_));
 sky130_fd_sc_hd__nand2_1 _07249_ (.A(net425),
    .B(net173),
    .Y(_01139_));
 sky130_fd_sc_hd__and4_1 _07250_ (.A(net185),
    .B(net429),
    .C(net165),
    .D(net620),
    .X(_01140_));
 sky130_fd_sc_hd__a22oi_1 _07251_ (.A1(net429),
    .A2(net165),
    .B1(net620),
    .B2(net185),
    .Y(_01141_));
 sky130_fd_sc_hd__nor2_1 _07252_ (.A(_01140_),
    .B(_01141_),
    .Y(_01142_));
 sky130_fd_sc_hd__xnor2_1 _07253_ (.A(_01139_),
    .B(_01142_),
    .Y(_01143_));
 sky130_fd_sc_hd__o21ba_1 _07254_ (.A1(_00985_),
    .A2(_00987_),
    .B1_N(_00986_),
    .X(_01144_));
 sky130_fd_sc_hd__and2b_1 _07255_ (.A_N(_01144_),
    .B(_01143_),
    .X(_01145_));
 sky130_fd_sc_hd__xnor2_1 _07256_ (.A(_01143_),
    .B(_01144_),
    .Y(_01146_));
 sky130_fd_sc_hd__and2_1 _07257_ (.A(_01138_),
    .B(_01146_),
    .X(_01147_));
 sky130_fd_sc_hd__xnor2_1 _07258_ (.A(_01138_),
    .B(_01146_),
    .Y(_01149_));
 sky130_fd_sc_hd__a21o_2 _07259_ (.A1(_01009_),
    .A2(_01011_),
    .B1(_01149_),
    .X(_01150_));
 sky130_fd_sc_hd__nand3_1 _07260_ (.A(_01009_),
    .B(_01011_),
    .C(_01149_),
    .Y(_01151_));
 sky130_fd_sc_hd__o211ai_4 _07261_ (.A1(_00991_),
    .A2(_00993_),
    .B1(_01150_),
    .C1(_01151_),
    .Y(_01152_));
 sky130_fd_sc_hd__a211o_1 _07262_ (.A1(_01150_),
    .A2(_01151_),
    .B1(_00991_),
    .C1(_00993_),
    .X(_01153_));
 sky130_fd_sc_hd__o21ba_1 _07263_ (.A1(_01003_),
    .A2(_01005_),
    .B1_N(_01004_),
    .X(_01154_));
 sky130_fd_sc_hd__o21ba_1 _07264_ (.A1(_01013_),
    .A2(_01015_),
    .B1_N(_01014_),
    .X(_01155_));
 sky130_fd_sc_hd__nand2_1 _07265_ (.A(net193),
    .B(net612),
    .Y(_01156_));
 sky130_fd_sc_hd__and4_1 _07266_ (.A(net210),
    .B(net201),
    .C(net596),
    .D(net589),
    .X(_01157_));
 sky130_fd_sc_hd__a22oi_1 _07267_ (.A1(net201),
    .A2(net596),
    .B1(net589),
    .B2(net210),
    .Y(_01158_));
 sky130_fd_sc_hd__nor2_1 _07268_ (.A(_01157_),
    .B(_01158_),
    .Y(_01160_));
 sky130_fd_sc_hd__xnor2_1 _07269_ (.A(_01156_),
    .B(_01160_),
    .Y(_01161_));
 sky130_fd_sc_hd__nand2b_1 _07270_ (.A_N(_01155_),
    .B(_01161_),
    .Y(_01162_));
 sky130_fd_sc_hd__xnor2_1 _07271_ (.A(_01155_),
    .B(_01161_),
    .Y(_01163_));
 sky130_fd_sc_hd__nand2b_1 _07272_ (.A_N(_01154_),
    .B(_01163_),
    .Y(_01164_));
 sky130_fd_sc_hd__xnor2_1 _07273_ (.A(_01154_),
    .B(_01163_),
    .Y(_01165_));
 sky130_fd_sc_hd__nand2_1 _07274_ (.A(net216),
    .B(net581),
    .Y(_01166_));
 sky130_fd_sc_hd__and4_1 _07275_ (.A(net238),
    .B(net230),
    .C(net575),
    .D(net570),
    .X(_01167_));
 sky130_fd_sc_hd__a22oi_1 _07276_ (.A1(net230),
    .A2(net575),
    .B1(net569),
    .B2(net238),
    .Y(_01168_));
 sky130_fd_sc_hd__nor2_1 _07277_ (.A(_01167_),
    .B(_01168_),
    .Y(_01169_));
 sky130_fd_sc_hd__xnor2_1 _07278_ (.A(_01166_),
    .B(_01169_),
    .Y(_01171_));
 sky130_fd_sc_hd__and2_1 _07279_ (.A(net257),
    .B(net562),
    .X(_01172_));
 sky130_fd_sc_hd__nand4_1 _07280_ (.A(net436),
    .B(net343),
    .C(net554),
    .D(net540),
    .Y(_01173_));
 sky130_fd_sc_hd__a22o_1 _07281_ (.A1(net343),
    .A2(net554),
    .B1(net540),
    .B2(net436),
    .X(_01174_));
 sky130_fd_sc_hd__nand3_1 _07282_ (.A(_01172_),
    .B(_01173_),
    .C(_01174_),
    .Y(_01175_));
 sky130_fd_sc_hd__a21o_1 _07283_ (.A1(_01173_),
    .A2(_01174_),
    .B1(_01172_),
    .X(_01176_));
 sky130_fd_sc_hd__o21bai_1 _07284_ (.A1(_01019_),
    .A2(_01021_),
    .B1_N(_01020_),
    .Y(_01177_));
 sky130_fd_sc_hd__nand3_1 _07285_ (.A(_01175_),
    .B(_01176_),
    .C(_01177_),
    .Y(_01178_));
 sky130_fd_sc_hd__a21o_1 _07286_ (.A1(_01175_),
    .A2(_01176_),
    .B1(_01177_),
    .X(_01179_));
 sky130_fd_sc_hd__nand3_1 _07287_ (.A(_01171_),
    .B(_01178_),
    .C(_01179_),
    .Y(_01180_));
 sky130_fd_sc_hd__a21o_1 _07288_ (.A1(_01178_),
    .A2(_01179_),
    .B1(_01171_),
    .X(_01182_));
 sky130_fd_sc_hd__a21bo_1 _07289_ (.A1(_01018_),
    .A2(_01026_),
    .B1_N(_01025_),
    .X(_01183_));
 sky130_fd_sc_hd__nand3_2 _07290_ (.A(_01180_),
    .B(_01182_),
    .C(_01183_),
    .Y(_01184_));
 sky130_fd_sc_hd__a21o_1 _07291_ (.A1(_01180_),
    .A2(_01182_),
    .B1(_01183_),
    .X(_01185_));
 sky130_fd_sc_hd__and3_1 _07292_ (.A(_01165_),
    .B(_01184_),
    .C(_01185_),
    .X(_01186_));
 sky130_fd_sc_hd__nand3_1 _07293_ (.A(_01165_),
    .B(_01184_),
    .C(_01185_),
    .Y(_01187_));
 sky130_fd_sc_hd__a21oi_1 _07294_ (.A1(_01184_),
    .A2(_01185_),
    .B1(_01165_),
    .Y(_01188_));
 sky130_fd_sc_hd__a211oi_1 _07295_ (.A1(_01031_),
    .A2(_01034_),
    .B1(_01186_),
    .C1(_01188_),
    .Y(_01189_));
 sky130_fd_sc_hd__a211o_1 _07296_ (.A1(_01031_),
    .A2(_01034_),
    .B1(_01186_),
    .C1(_01188_),
    .X(_01190_));
 sky130_fd_sc_hd__o211ai_2 _07297_ (.A1(_01186_),
    .A2(_01188_),
    .B1(_01031_),
    .C1(_01034_),
    .Y(_01191_));
 sky130_fd_sc_hd__and4_1 _07298_ (.A(_01152_),
    .B(_01153_),
    .C(_01190_),
    .D(_01191_),
    .X(_01193_));
 sky130_fd_sc_hd__a22oi_2 _07299_ (.A1(_01152_),
    .A2(_01153_),
    .B1(_01190_),
    .B2(_01191_),
    .Y(_01194_));
 sky130_fd_sc_hd__a211o_1 _07300_ (.A1(_01036_),
    .A2(_01038_),
    .B1(_01193_),
    .C1(_01194_),
    .X(_01195_));
 sky130_fd_sc_hd__o211ai_1 _07301_ (.A1(_01193_),
    .A2(_01194_),
    .B1(_01036_),
    .C1(_01038_),
    .Y(_01196_));
 sky130_fd_sc_hd__or4bb_4 _07302_ (.A(_01131_),
    .B(_01132_),
    .C_N(_01195_),
    .D_N(_01196_),
    .X(_01197_));
 sky130_fd_sc_hd__a2bb2o_1 _07303_ (.A1_N(_01131_),
    .A2_N(_01132_),
    .B1(_01195_),
    .B2(_01196_),
    .X(_01198_));
 sky130_fd_sc_hd__o211ai_4 _07304_ (.A1(_01041_),
    .A2(net139),
    .B1(_01197_),
    .C1(_01198_),
    .Y(_01199_));
 sky130_fd_sc_hd__a211o_1 _07305_ (.A1(_01197_),
    .A2(_01198_),
    .B1(_01041_),
    .C1(_01043_),
    .X(_01200_));
 sky130_fd_sc_hd__nand4_2 _07306_ (.A(_01092_),
    .B(_01094_),
    .C(_01199_),
    .D(_01200_),
    .Y(_01201_));
 sky130_fd_sc_hd__a22o_1 _07307_ (.A1(_01092_),
    .A2(_01094_),
    .B1(_01199_),
    .B2(_01200_),
    .X(_01202_));
 sky130_fd_sc_hd__o211a_1 _07308_ (.A1(_01045_),
    .A2(_01047_),
    .B1(_01201_),
    .C1(_01202_),
    .X(_01204_));
 sky130_fd_sc_hd__a211oi_1 _07309_ (.A1(_01201_),
    .A2(_01202_),
    .B1(_01045_),
    .C1(_01047_),
    .Y(_01205_));
 sky130_fd_sc_hd__a211oi_2 _07310_ (.A1(_00937_),
    .A2(_00939_),
    .B1(_01204_),
    .C1(_01205_),
    .Y(_01206_));
 sky130_fd_sc_hd__o211a_1 _07311_ (.A1(_01204_),
    .A2(_01205_),
    .B1(_00937_),
    .C1(_00939_),
    .X(_01207_));
 sky130_fd_sc_hd__a211oi_2 _07312_ (.A1(_01051_),
    .A2(_01053_),
    .B1(_01206_),
    .C1(_01207_),
    .Y(_01208_));
 sky130_fd_sc_hd__o211a_1 _07313_ (.A1(_01206_),
    .A2(_01207_),
    .B1(_01051_),
    .C1(_01053_),
    .X(_01209_));
 sky130_fd_sc_hd__o21ba_1 _07314_ (.A1(_01208_),
    .A2(_01209_),
    .B1_N(_01055_),
    .X(_01210_));
 sky130_fd_sc_hd__or3b_1 _07315_ (.A(_01208_),
    .B(_01209_),
    .C_N(_01055_),
    .X(_01211_));
 sky130_fd_sc_hd__inv_2 _07316_ (.A(_01211_),
    .Y(_01212_));
 sky130_fd_sc_hd__nor2_1 _07317_ (.A(_01210_),
    .B(_01212_),
    .Y(_01213_));
 sky130_fd_sc_hd__nor2_1 _07318_ (.A(_01058_),
    .B(_01064_),
    .Y(_01215_));
 sky130_fd_sc_hd__xnor2_1 _07319_ (.A(_01213_),
    .B(_01215_),
    .Y(net84));
 sky130_fd_sc_hd__o21ba_1 _07320_ (.A1(_01058_),
    .A2(_01212_),
    .B1_N(_01210_),
    .X(_01216_));
 sky130_fd_sc_hd__a21oi_2 _07321_ (.A1(_01064_),
    .A2(_01213_),
    .B1(_01216_),
    .Y(_01217_));
 sky130_fd_sc_hd__and2b_1 _07322_ (.A_N(_01091_),
    .B(_01094_),
    .X(_01218_));
 sky130_fd_sc_hd__a22o_1 _07323_ (.A1(net603),
    .A2(net282),
    .B1(net273),
    .B2(net631),
    .X(_01219_));
 sky130_fd_sc_hd__and4_1 _07324_ (.A(net603),
    .B(net628),
    .C(net282),
    .D(net273),
    .X(_01220_));
 sky130_fd_sc_hd__nand4_1 _07325_ (.A(net603),
    .B(net631),
    .C(net282),
    .D(net273),
    .Y(_01221_));
 sky130_fd_sc_hd__nor2_1 _07326_ (.A(_01069_),
    .B(_01073_),
    .Y(_01222_));
 sky130_fd_sc_hd__nor2_1 _07327_ (.A(_01095_),
    .B(_01097_),
    .Y(_01223_));
 sky130_fd_sc_hd__and4_1 _07328_ (.A(net488),
    .B(net497),
    .C(net310),
    .D(net296),
    .X(_01225_));
 sky130_fd_sc_hd__a22oi_1 _07329_ (.A1(net489),
    .A2(net310),
    .B1(net296),
    .B2(net497),
    .Y(_01226_));
 sky130_fd_sc_hd__nor2_1 _07330_ (.A(_01225_),
    .B(_01226_),
    .Y(_01227_));
 sky130_fd_sc_hd__nand2_1 _07331_ (.A(net517),
    .B(net288),
    .Y(_01228_));
 sky130_fd_sc_hd__xnor2_1 _07332_ (.A(_01227_),
    .B(_01228_),
    .Y(_01229_));
 sky130_fd_sc_hd__nand2b_1 _07333_ (.A_N(_01223_),
    .B(_01229_),
    .Y(_01230_));
 sky130_fd_sc_hd__xnor2_1 _07334_ (.A(_01223_),
    .B(_01229_),
    .Y(_01231_));
 sky130_fd_sc_hd__nand2b_1 _07335_ (.A_N(_01222_),
    .B(_01231_),
    .Y(_01232_));
 sky130_fd_sc_hd__xnor2_1 _07336_ (.A(_01222_),
    .B(_01231_),
    .Y(_01233_));
 sky130_fd_sc_hd__o21a_1 _07337_ (.A1(_01107_),
    .A2(_01109_),
    .B1(_01233_),
    .X(_01234_));
 sky130_fd_sc_hd__o21ai_1 _07338_ (.A1(_01107_),
    .A2(_01109_),
    .B1(_01233_),
    .Y(_01236_));
 sky130_fd_sc_hd__nor3_1 _07339_ (.A(_01107_),
    .B(_01109_),
    .C(_01233_),
    .Y(_01237_));
 sky130_fd_sc_hd__a211o_2 _07340_ (.A1(_01075_),
    .A2(_01077_),
    .B1(_01234_),
    .C1(_01237_),
    .X(_01238_));
 sky130_fd_sc_hd__o211ai_2 _07341_ (.A1(_01234_),
    .A2(_01237_),
    .B1(_01075_),
    .C1(_01077_),
    .Y(_01239_));
 sky130_fd_sc_hd__o211ai_4 _07342_ (.A1(_01079_),
    .A2(_01081_),
    .B1(_01238_),
    .C1(_01239_),
    .Y(_01240_));
 sky130_fd_sc_hd__a211o_1 _07343_ (.A1(_01238_),
    .A2(_01239_),
    .B1(_01079_),
    .C1(_01081_),
    .X(_01241_));
 sky130_fd_sc_hd__nand4_2 _07344_ (.A(_01219_),
    .B(_01221_),
    .C(_01240_),
    .D(_01241_),
    .Y(_01242_));
 sky130_fd_sc_hd__a22o_1 _07345_ (.A1(_01219_),
    .A2(_01221_),
    .B1(_01240_),
    .B2(_01241_),
    .X(_01243_));
 sky130_fd_sc_hd__o211a_1 _07346_ (.A1(_01129_),
    .A2(_01131_),
    .B1(_01242_),
    .C1(_01243_),
    .X(_01244_));
 sky130_fd_sc_hd__inv_2 _07347_ (.A(_01244_),
    .Y(_01245_));
 sky130_fd_sc_hd__a211oi_1 _07348_ (.A1(_01242_),
    .A2(_01243_),
    .B1(_01129_),
    .C1(_01131_),
    .Y(_01247_));
 sky130_fd_sc_hd__a211o_1 _07349_ (.A1(_01085_),
    .A2(_01088_),
    .B1(_01244_),
    .C1(_01247_),
    .X(_01248_));
 sky130_fd_sc_hd__o211ai_2 _07350_ (.A1(_01244_),
    .A2(_01247_),
    .B1(_01085_),
    .C1(_01088_),
    .Y(_01249_));
 sky130_fd_sc_hd__nand2_1 _07351_ (.A(net482),
    .B(net48),
    .Y(_01250_));
 sky130_fd_sc_hd__and4_1 _07352_ (.A(net474),
    .B(net461),
    .C(net330),
    .D(net323),
    .X(_01251_));
 sky130_fd_sc_hd__a22oi_1 _07353_ (.A1(net461),
    .A2(net330),
    .B1(net323),
    .B2(net474),
    .Y(_01252_));
 sky130_fd_sc_hd__nor2_1 _07354_ (.A(_01251_),
    .B(_01252_),
    .Y(_01253_));
 sky130_fd_sc_hd__xnor2_1 _07355_ (.A(_01250_),
    .B(_01253_),
    .Y(_01254_));
 sky130_fd_sc_hd__nand2_1 _07356_ (.A(net455),
    .B(net339),
    .Y(_01255_));
 sky130_fd_sc_hd__and4_1 _07357_ (.A(net549),
    .B(net448),
    .C(net361),
    .D(net353),
    .X(_01256_));
 sky130_fd_sc_hd__a22oi_1 _07358_ (.A1(net549),
    .A2(net361),
    .B1(net353),
    .B2(net448),
    .Y(_01258_));
 sky130_fd_sc_hd__nor2_1 _07359_ (.A(_01256_),
    .B(_01258_),
    .Y(_01259_));
 sky130_fd_sc_hd__xnor2_1 _07360_ (.A(_01255_),
    .B(_01259_),
    .Y(_01260_));
 sky130_fd_sc_hd__o21ba_1 _07361_ (.A1(_01100_),
    .A2(_01102_),
    .B1_N(_01101_),
    .X(_01261_));
 sky130_fd_sc_hd__and2b_1 _07362_ (.A_N(_01261_),
    .B(_01260_),
    .X(_01262_));
 sky130_fd_sc_hd__xnor2_1 _07363_ (.A(_01260_),
    .B(_01261_),
    .Y(_01263_));
 sky130_fd_sc_hd__and2_1 _07364_ (.A(_01254_),
    .B(_01263_),
    .X(_01264_));
 sky130_fd_sc_hd__nor2_1 _07365_ (.A(_01254_),
    .B(_01263_),
    .Y(_01265_));
 sky130_fd_sc_hd__or2_1 _07366_ (.A(_01264_),
    .B(_01265_),
    .X(_01266_));
 sky130_fd_sc_hd__a31o_1 _07367_ (.A1(net549),
    .A2(net369),
    .A3(_01118_),
    .B1(_01116_),
    .X(_01267_));
 sky130_fd_sc_hd__o21ba_1 _07368_ (.A1(_01133_),
    .A2(_01135_),
    .B1_N(_01134_),
    .X(_01269_));
 sky130_fd_sc_hd__a22oi_1 _07369_ (.A1(net301),
    .A2(net392),
    .B1(net376),
    .B2(net386),
    .Y(_01270_));
 sky130_fd_sc_hd__and4_1 _07370_ (.A(net386),
    .B(net301),
    .C(net392),
    .D(net377),
    .X(_01271_));
 sky130_fd_sc_hd__nor2_1 _07371_ (.A(_01270_),
    .B(_01271_),
    .Y(_01272_));
 sky130_fd_sc_hd__nand2_1 _07372_ (.A(net468),
    .B(net369),
    .Y(_01273_));
 sky130_fd_sc_hd__xnor2_1 _07373_ (.A(_01272_),
    .B(_01273_),
    .Y(_01274_));
 sky130_fd_sc_hd__nand2b_1 _07374_ (.A_N(_01269_),
    .B(_01274_),
    .Y(_01275_));
 sky130_fd_sc_hd__xnor2_1 _07375_ (.A(_01269_),
    .B(_01274_),
    .Y(_01276_));
 sky130_fd_sc_hd__nand2_1 _07376_ (.A(_01267_),
    .B(_01276_),
    .Y(_01277_));
 sky130_fd_sc_hd__xnor2_1 _07377_ (.A(_01267_),
    .B(_01276_),
    .Y(_01278_));
 sky130_fd_sc_hd__a21oi_1 _07378_ (.A1(_01120_),
    .A2(_01122_),
    .B1(_01278_),
    .Y(_01279_));
 sky130_fd_sc_hd__and3_1 _07379_ (.A(_01120_),
    .B(_01122_),
    .C(_01278_),
    .X(_01280_));
 sky130_fd_sc_hd__nor3_1 _07380_ (.A(_01266_),
    .B(_01279_),
    .C(_01280_),
    .Y(_01281_));
 sky130_fd_sc_hd__o21a_1 _07381_ (.A1(_01279_),
    .A2(_01280_),
    .B1(_01266_),
    .X(_01282_));
 sky130_fd_sc_hd__a211oi_2 _07382_ (.A1(_01150_),
    .A2(_01152_),
    .B1(_01281_),
    .C1(_01282_),
    .Y(_01283_));
 sky130_fd_sc_hd__o211a_1 _07383_ (.A1(_01281_),
    .A2(_01282_),
    .B1(_01150_),
    .C1(_01152_),
    .X(_01284_));
 sky130_fd_sc_hd__a211oi_2 _07384_ (.A1(_01124_),
    .A2(_01127_),
    .B1(_01283_),
    .C1(_01284_),
    .Y(_01285_));
 sky130_fd_sc_hd__o211a_1 _07385_ (.A1(_01283_),
    .A2(_01284_),
    .B1(_01124_),
    .C1(_01127_),
    .X(_01286_));
 sky130_fd_sc_hd__nand2_1 _07386_ (.A(net225),
    .B(net401),
    .Y(_01287_));
 sky130_fd_sc_hd__and4_1 _07387_ (.A(net416),
    .B(net408),
    .C(net180),
    .D(net173),
    .X(_01288_));
 sky130_fd_sc_hd__a22oi_1 _07388_ (.A1(net408),
    .A2(net180),
    .B1(net173),
    .B2(net416),
    .Y(_01290_));
 sky130_fd_sc_hd__nor2_1 _07389_ (.A(_01288_),
    .B(_01290_),
    .Y(_01291_));
 sky130_fd_sc_hd__xnor2_1 _07390_ (.A(_01287_),
    .B(_01291_),
    .Y(_01292_));
 sky130_fd_sc_hd__nand2_1 _07391_ (.A(net422),
    .B(net165),
    .Y(_01293_));
 sky130_fd_sc_hd__and4_1 _07392_ (.A(net183),
    .B(net427),
    .C(net620),
    .D(net612),
    .X(_01294_));
 sky130_fd_sc_hd__a22o_1 _07393_ (.A1(net427),
    .A2(net620),
    .B1(net612),
    .B2(net183),
    .X(_01295_));
 sky130_fd_sc_hd__and2b_1 _07394_ (.A_N(_01294_),
    .B(_01295_),
    .X(_01296_));
 sky130_fd_sc_hd__xnor2_1 _07395_ (.A(_01293_),
    .B(_01296_),
    .Y(_01297_));
 sky130_fd_sc_hd__o21ba_1 _07396_ (.A1(_01139_),
    .A2(_01141_),
    .B1_N(_01140_),
    .X(_01298_));
 sky130_fd_sc_hd__and2b_1 _07397_ (.A_N(_01298_),
    .B(_01297_),
    .X(_01299_));
 sky130_fd_sc_hd__xnor2_1 _07398_ (.A(_01297_),
    .B(_01298_),
    .Y(_01301_));
 sky130_fd_sc_hd__and2_1 _07399_ (.A(_01292_),
    .B(_01301_),
    .X(_01302_));
 sky130_fd_sc_hd__xnor2_1 _07400_ (.A(_01292_),
    .B(_01301_),
    .Y(_01303_));
 sky130_fd_sc_hd__a21oi_1 _07401_ (.A1(_01162_),
    .A2(_01164_),
    .B1(_01303_),
    .Y(_01304_));
 sky130_fd_sc_hd__a21o_1 _07402_ (.A1(_01162_),
    .A2(_01164_),
    .B1(_01303_),
    .X(_01305_));
 sky130_fd_sc_hd__nand3_1 _07403_ (.A(_01162_),
    .B(_01164_),
    .C(_01303_),
    .Y(_01306_));
 sky130_fd_sc_hd__o211a_1 _07404_ (.A1(_01145_),
    .A2(_01147_),
    .B1(_01305_),
    .C1(_01306_),
    .X(_01307_));
 sky130_fd_sc_hd__a211oi_1 _07405_ (.A1(_01305_),
    .A2(_01306_),
    .B1(_01145_),
    .C1(_01147_),
    .Y(_01308_));
 sky130_fd_sc_hd__a31o_1 _07406_ (.A1(net193),
    .A2(net612),
    .A3(_01160_),
    .B1(_01157_),
    .X(_01309_));
 sky130_fd_sc_hd__o21bai_1 _07407_ (.A1(_01166_),
    .A2(_01168_),
    .B1_N(_01167_),
    .Y(_01310_));
 sky130_fd_sc_hd__nand2_1 _07408_ (.A(net193),
    .B(net596),
    .Y(_01312_));
 sky130_fd_sc_hd__nand4_1 _07409_ (.A(net210),
    .B(net201),
    .C(net589),
    .D(net581),
    .Y(_01313_));
 sky130_fd_sc_hd__a22o_1 _07410_ (.A1(net201),
    .A2(net589),
    .B1(net581),
    .B2(net210),
    .X(_01314_));
 sky130_fd_sc_hd__nand3b_1 _07411_ (.A_N(_01312_),
    .B(_01313_),
    .C(_01314_),
    .Y(_01315_));
 sky130_fd_sc_hd__a21bo_1 _07412_ (.A1(_01313_),
    .A2(_01314_),
    .B1_N(_01312_),
    .X(_01316_));
 sky130_fd_sc_hd__and3_1 _07413_ (.A(_01310_),
    .B(_01315_),
    .C(_01316_),
    .X(_01317_));
 sky130_fd_sc_hd__a21o_1 _07414_ (.A1(_01315_),
    .A2(_01316_),
    .B1(_01310_),
    .X(_01318_));
 sky130_fd_sc_hd__and2b_1 _07415_ (.A_N(_01317_),
    .B(_01318_),
    .X(_01319_));
 sky130_fd_sc_hd__xor2_1 _07416_ (.A(_01309_),
    .B(_01319_),
    .X(_01320_));
 sky130_fd_sc_hd__nand2_1 _07417_ (.A(net216),
    .B(net575),
    .Y(_01321_));
 sky130_fd_sc_hd__and4_1 _07418_ (.A(net237),
    .B(net230),
    .C(net568),
    .D(net562),
    .X(_01323_));
 sky130_fd_sc_hd__a22oi_1 _07419_ (.A1(net230),
    .A2(net568),
    .B1(net562),
    .B2(net237),
    .Y(_01324_));
 sky130_fd_sc_hd__nor2_1 _07420_ (.A(_01323_),
    .B(_01324_),
    .Y(_01325_));
 sky130_fd_sc_hd__xnor2_1 _07421_ (.A(_01321_),
    .B(_01325_),
    .Y(_01326_));
 sky130_fd_sc_hd__nand2_1 _07422_ (.A(net257),
    .B(net554),
    .Y(_01327_));
 sky130_fd_sc_hd__and4_1 _07423_ (.A(net436),
    .B(net344),
    .C(net540),
    .D(net534),
    .X(_01328_));
 sky130_fd_sc_hd__a22oi_2 _07424_ (.A1(net344),
    .A2(net540),
    .B1(net534),
    .B2(net436),
    .Y(_01329_));
 sky130_fd_sc_hd__or3_1 _07425_ (.A(_01327_),
    .B(_01328_),
    .C(_01329_),
    .X(_01330_));
 sky130_fd_sc_hd__o21ai_1 _07426_ (.A1(_01328_),
    .A2(_01329_),
    .B1(_01327_),
    .Y(_01331_));
 sky130_fd_sc_hd__a21bo_1 _07427_ (.A1(_01172_),
    .A2(_01174_),
    .B1_N(_01173_),
    .X(_01332_));
 sky130_fd_sc_hd__nand3_1 _07428_ (.A(_01330_),
    .B(_01331_),
    .C(_01332_),
    .Y(_01334_));
 sky130_fd_sc_hd__a21o_1 _07429_ (.A1(_01330_),
    .A2(_01331_),
    .B1(_01332_),
    .X(_01335_));
 sky130_fd_sc_hd__nand3_1 _07430_ (.A(_01326_),
    .B(_01334_),
    .C(_01335_),
    .Y(_01336_));
 sky130_fd_sc_hd__a21o_1 _07431_ (.A1(_01334_),
    .A2(_01335_),
    .B1(_01326_),
    .X(_01337_));
 sky130_fd_sc_hd__a21bo_1 _07432_ (.A1(_01171_),
    .A2(_01179_),
    .B1_N(_01178_),
    .X(_01338_));
 sky130_fd_sc_hd__nand3_2 _07433_ (.A(_01336_),
    .B(_01337_),
    .C(_01338_),
    .Y(_01339_));
 sky130_fd_sc_hd__a21o_1 _07434_ (.A1(_01336_),
    .A2(_01337_),
    .B1(_01338_),
    .X(_01340_));
 sky130_fd_sc_hd__and3_1 _07435_ (.A(_01320_),
    .B(_01339_),
    .C(_01340_),
    .X(_01341_));
 sky130_fd_sc_hd__nand3_2 _07436_ (.A(_01320_),
    .B(_01339_),
    .C(_01340_),
    .Y(_01342_));
 sky130_fd_sc_hd__a21oi_1 _07437_ (.A1(_01339_),
    .A2(_01340_),
    .B1(_01320_),
    .Y(_01343_));
 sky130_fd_sc_hd__a211o_1 _07438_ (.A1(_01184_),
    .A2(_01187_),
    .B1(_01341_),
    .C1(_01343_),
    .X(_01345_));
 sky130_fd_sc_hd__o211ai_1 _07439_ (.A1(_01341_),
    .A2(_01343_),
    .B1(_01184_),
    .C1(_01187_),
    .Y(_01346_));
 sky130_fd_sc_hd__or4bb_2 _07440_ (.A(_01307_),
    .B(_01308_),
    .C_N(_01345_),
    .D_N(_01346_),
    .X(_01347_));
 sky130_fd_sc_hd__a2bb2o_1 _07441_ (.A1_N(_01307_),
    .A2_N(_01308_),
    .B1(_01345_),
    .B2(_01346_),
    .X(_01348_));
 sky130_fd_sc_hd__o211a_1 _07442_ (.A1(_01189_),
    .A2(_01193_),
    .B1(_01347_),
    .C1(_01348_),
    .X(_01349_));
 sky130_fd_sc_hd__a211oi_1 _07443_ (.A1(_01347_),
    .A2(_01348_),
    .B1(_01189_),
    .C1(_01193_),
    .Y(_01350_));
 sky130_fd_sc_hd__nor4_1 _07444_ (.A(_01285_),
    .B(_01286_),
    .C(_01349_),
    .D(_01350_),
    .Y(_01351_));
 sky130_fd_sc_hd__o22a_1 _07445_ (.A1(_01285_),
    .A2(_01286_),
    .B1(_01349_),
    .B2(_01350_),
    .X(_01352_));
 sky130_fd_sc_hd__a211oi_1 _07446_ (.A1(_01195_),
    .A2(_01197_),
    .B1(net138),
    .C1(_01352_),
    .Y(_01353_));
 sky130_fd_sc_hd__a211o_1 _07447_ (.A1(_01195_),
    .A2(_01197_),
    .B1(net138),
    .C1(_01352_),
    .X(_01354_));
 sky130_fd_sc_hd__o211ai_1 _07448_ (.A1(net138),
    .A2(_01352_),
    .B1(_01195_),
    .C1(_01197_),
    .Y(_01356_));
 sky130_fd_sc_hd__and4_1 _07449_ (.A(_01248_),
    .B(_01249_),
    .C(_01354_),
    .D(_01356_),
    .X(_01357_));
 sky130_fd_sc_hd__a22oi_2 _07450_ (.A1(_01248_),
    .A2(_01249_),
    .B1(_01354_),
    .B2(_01356_),
    .Y(_01358_));
 sky130_fd_sc_hd__a211oi_1 _07451_ (.A1(_01199_),
    .A2(_01201_),
    .B1(_01357_),
    .C1(_01358_),
    .Y(_01359_));
 sky130_fd_sc_hd__a211o_1 _07452_ (.A1(_01199_),
    .A2(_01201_),
    .B1(_01357_),
    .C1(_01358_),
    .X(_01360_));
 sky130_fd_sc_hd__o211a_1 _07453_ (.A1(_01357_),
    .A2(_01358_),
    .B1(_01199_),
    .C1(_01201_),
    .X(_01361_));
 sky130_fd_sc_hd__or3_2 _07454_ (.A(_01218_),
    .B(_01359_),
    .C(_01361_),
    .X(_01362_));
 sky130_fd_sc_hd__o21ai_1 _07455_ (.A1(_01359_),
    .A2(_01361_),
    .B1(_01218_),
    .Y(_01363_));
 sky130_fd_sc_hd__o211a_1 _07456_ (.A1(_01204_),
    .A2(_01206_),
    .B1(_01362_),
    .C1(_01363_),
    .X(_01364_));
 sky130_fd_sc_hd__a211oi_1 _07457_ (.A1(_01362_),
    .A2(_01363_),
    .B1(_01204_),
    .C1(_01206_),
    .Y(_01365_));
 sky130_fd_sc_hd__nor3b_1 _07458_ (.A(_01364_),
    .B(_01365_),
    .C_N(_01208_),
    .Y(_01367_));
 sky130_fd_sc_hd__o21ba_1 _07459_ (.A1(_01364_),
    .A2(_01365_),
    .B1_N(_01208_),
    .X(_01368_));
 sky130_fd_sc_hd__or2_1 _07460_ (.A(_01367_),
    .B(_01368_),
    .X(_01369_));
 sky130_fd_sc_hd__xor2_1 _07461_ (.A(_01217_),
    .B(_01369_),
    .X(net85));
 sky130_fd_sc_hd__and4_1 _07462_ (.A(net520),
    .B(net602),
    .C(net282),
    .D(net273),
    .X(_01370_));
 sky130_fd_sc_hd__a22oi_1 _07463_ (.A1(net520),
    .A2(net282),
    .B1(net273),
    .B2(net602),
    .Y(_01371_));
 sky130_fd_sc_hd__nor2_1 _07464_ (.A(_01370_),
    .B(_01371_),
    .Y(_01372_));
 sky130_fd_sc_hd__nand2_1 _07465_ (.A(net628),
    .B(net264),
    .Y(_01373_));
 sky130_fd_sc_hd__xnor2_1 _07466_ (.A(_01372_),
    .B(_01373_),
    .Y(_01374_));
 sky130_fd_sc_hd__nand2_1 _07467_ (.A(_01220_),
    .B(_01374_),
    .Y(_01375_));
 sky130_fd_sc_hd__or2_1 _07468_ (.A(_01220_),
    .B(_01374_),
    .X(_01377_));
 sky130_fd_sc_hd__nand2_1 _07469_ (.A(_01375_),
    .B(_01377_),
    .Y(_01378_));
 sky130_fd_sc_hd__o21ba_1 _07470_ (.A1(_01226_),
    .A2(_01228_),
    .B1_N(_01225_),
    .X(_01379_));
 sky130_fd_sc_hd__o21ba_1 _07471_ (.A1(_01250_),
    .A2(_01252_),
    .B1_N(_01251_),
    .X(_01380_));
 sky130_fd_sc_hd__and4_1 _07472_ (.A(net482),
    .B(net489),
    .C(net308),
    .D(net50),
    .X(_01381_));
 sky130_fd_sc_hd__a22oi_1 _07473_ (.A1(net482),
    .A2(net310),
    .B1(net50),
    .B2(net489),
    .Y(_01382_));
 sky130_fd_sc_hd__nor2_1 _07474_ (.A(_01381_),
    .B(_01382_),
    .Y(_01383_));
 sky130_fd_sc_hd__nand2_1 _07475_ (.A(net497),
    .B(net288),
    .Y(_01384_));
 sky130_fd_sc_hd__xnor2_1 _07476_ (.A(_01383_),
    .B(_01384_),
    .Y(_01385_));
 sky130_fd_sc_hd__nand2b_1 _07477_ (.A_N(_01380_),
    .B(_01385_),
    .Y(_01386_));
 sky130_fd_sc_hd__xnor2_1 _07478_ (.A(_01380_),
    .B(_01385_),
    .Y(_01388_));
 sky130_fd_sc_hd__nand2b_1 _07479_ (.A_N(_01379_),
    .B(_01388_),
    .Y(_01389_));
 sky130_fd_sc_hd__xnor2_1 _07480_ (.A(_01379_),
    .B(_01388_),
    .Y(_01390_));
 sky130_fd_sc_hd__o21a_1 _07481_ (.A1(_01262_),
    .A2(_01264_),
    .B1(_01390_),
    .X(_01391_));
 sky130_fd_sc_hd__nor3_1 _07482_ (.A(_01262_),
    .B(_01264_),
    .C(_01390_),
    .Y(_01392_));
 sky130_fd_sc_hd__a211oi_2 _07483_ (.A1(_01230_),
    .A2(_01232_),
    .B1(_01391_),
    .C1(_01392_),
    .Y(_01393_));
 sky130_fd_sc_hd__o211a_1 _07484_ (.A1(_01391_),
    .A2(_01392_),
    .B1(_01230_),
    .C1(_01232_),
    .X(_01394_));
 sky130_fd_sc_hd__a211oi_1 _07485_ (.A1(_01236_),
    .A2(_01238_),
    .B1(_01393_),
    .C1(_01394_),
    .Y(_01395_));
 sky130_fd_sc_hd__a211o_1 _07486_ (.A1(_01236_),
    .A2(_01238_),
    .B1(_01393_),
    .C1(_01394_),
    .X(_01396_));
 sky130_fd_sc_hd__o211a_1 _07487_ (.A1(_01393_),
    .A2(_01394_),
    .B1(_01236_),
    .C1(_01238_),
    .X(_01397_));
 sky130_fd_sc_hd__or3_1 _07488_ (.A(_01378_),
    .B(_01395_),
    .C(_01397_),
    .X(_01399_));
 sky130_fd_sc_hd__o21ai_1 _07489_ (.A1(_01395_),
    .A2(_01397_),
    .B1(_01378_),
    .Y(_01400_));
 sky130_fd_sc_hd__o211a_1 _07490_ (.A1(_01283_),
    .A2(_01285_),
    .B1(_01399_),
    .C1(_01400_),
    .X(_01401_));
 sky130_fd_sc_hd__a211oi_1 _07491_ (.A1(_01399_),
    .A2(_01400_),
    .B1(_01283_),
    .C1(_01285_),
    .Y(_01402_));
 sky130_fd_sc_hd__a211oi_2 _07492_ (.A1(_01240_),
    .A2(_01242_),
    .B1(_01401_),
    .C1(_01402_),
    .Y(_01403_));
 sky130_fd_sc_hd__o211a_1 _07493_ (.A1(_01401_),
    .A2(_01402_),
    .B1(_01240_),
    .C1(_01242_),
    .X(_01404_));
 sky130_fd_sc_hd__nor2_1 _07494_ (.A(_01279_),
    .B(_01281_),
    .Y(_01405_));
 sky130_fd_sc_hd__and4_1 _07495_ (.A(net459),
    .B(net450),
    .C(net331),
    .D(net324),
    .X(_01406_));
 sky130_fd_sc_hd__a22o_1 _07496_ (.A1(net450),
    .A2(net331),
    .B1(net324),
    .B2(net459),
    .X(_01407_));
 sky130_fd_sc_hd__and2b_1 _07497_ (.A_N(_01406_),
    .B(_01407_),
    .X(_01408_));
 sky130_fd_sc_hd__nand2_1 _07498_ (.A(net474),
    .B(net316),
    .Y(_01410_));
 sky130_fd_sc_hd__xnor2_1 _07499_ (.A(_01408_),
    .B(_01410_),
    .Y(_01411_));
 sky130_fd_sc_hd__nand2_1 _07500_ (.A(net443),
    .B(net339),
    .Y(_01412_));
 sky130_fd_sc_hd__and4_1 _07501_ (.A(net544),
    .B(net468),
    .C(net42),
    .D(net43),
    .X(_01413_));
 sky130_fd_sc_hd__a22oi_2 _07502_ (.A1(net468),
    .A2(net362),
    .B1(net354),
    .B2(net544),
    .Y(_01414_));
 sky130_fd_sc_hd__or3_1 _07503_ (.A(_01412_),
    .B(_01413_),
    .C(_01414_),
    .X(_01415_));
 sky130_fd_sc_hd__o21ai_1 _07504_ (.A1(_01413_),
    .A2(_01414_),
    .B1(_01412_),
    .Y(_01416_));
 sky130_fd_sc_hd__o21bai_1 _07505_ (.A1(_01255_),
    .A2(_01258_),
    .B1_N(_01256_),
    .Y(_01417_));
 sky130_fd_sc_hd__and3_1 _07506_ (.A(_01415_),
    .B(_01416_),
    .C(_01417_),
    .X(_01418_));
 sky130_fd_sc_hd__a21o_1 _07507_ (.A1(_01415_),
    .A2(_01416_),
    .B1(_01417_),
    .X(_01419_));
 sky130_fd_sc_hd__and2b_1 _07508_ (.A_N(_01418_),
    .B(_01419_),
    .X(_01421_));
 sky130_fd_sc_hd__xnor2_1 _07509_ (.A(_01411_),
    .B(_01421_),
    .Y(_01422_));
 sky130_fd_sc_hd__a31o_1 _07510_ (.A1(net468),
    .A2(net369),
    .A3(_01272_),
    .B1(_01271_),
    .X(_01423_));
 sky130_fd_sc_hd__o21bai_1 _07511_ (.A1(_01287_),
    .A2(_01290_),
    .B1_N(_01288_),
    .Y(_01424_));
 sky130_fd_sc_hd__nand4_1 _07512_ (.A(net301),
    .B(net225),
    .C(net393),
    .D(net377),
    .Y(_01425_));
 sky130_fd_sc_hd__a22o_1 _07513_ (.A1(net225),
    .A2(net393),
    .B1(net377),
    .B2(net301),
    .X(_01426_));
 sky130_fd_sc_hd__a22o_1 _07514_ (.A1(net386),
    .A2(net369),
    .B1(_01425_),
    .B2(_01426_),
    .X(_01427_));
 sky130_fd_sc_hd__nand4_1 _07515_ (.A(net386),
    .B(net372),
    .C(_01425_),
    .D(_01426_),
    .Y(_01428_));
 sky130_fd_sc_hd__nand3_1 _07516_ (.A(_01424_),
    .B(_01427_),
    .C(_01428_),
    .Y(_01429_));
 sky130_fd_sc_hd__a21o_1 _07517_ (.A1(_01427_),
    .A2(_01428_),
    .B1(_01424_),
    .X(_01430_));
 sky130_fd_sc_hd__and3_1 _07518_ (.A(_01423_),
    .B(_01429_),
    .C(_01430_),
    .X(_01432_));
 sky130_fd_sc_hd__a21oi_1 _07519_ (.A1(_01429_),
    .A2(_01430_),
    .B1(_01423_),
    .Y(_01433_));
 sky130_fd_sc_hd__or2_1 _07520_ (.A(_01432_),
    .B(_01433_),
    .X(_01434_));
 sky130_fd_sc_hd__a21oi_1 _07521_ (.A1(_01275_),
    .A2(_01277_),
    .B1(_01434_),
    .Y(_01435_));
 sky130_fd_sc_hd__a21o_1 _07522_ (.A1(_01275_),
    .A2(_01277_),
    .B1(_01434_),
    .X(_01436_));
 sky130_fd_sc_hd__and3_1 _07523_ (.A(_01275_),
    .B(_01277_),
    .C(_01434_),
    .X(_01437_));
 sky130_fd_sc_hd__or3_1 _07524_ (.A(_01422_),
    .B(_01435_),
    .C(_01437_),
    .X(_01438_));
 sky130_fd_sc_hd__o21ai_1 _07525_ (.A1(_01435_),
    .A2(_01437_),
    .B1(_01422_),
    .Y(_01439_));
 sky130_fd_sc_hd__o211a_1 _07526_ (.A1(_01304_),
    .A2(_01307_),
    .B1(_01438_),
    .C1(_01439_),
    .X(_01440_));
 sky130_fd_sc_hd__a211oi_1 _07527_ (.A1(_01438_),
    .A2(_01439_),
    .B1(_01304_),
    .C1(_01307_),
    .Y(_01441_));
 sky130_fd_sc_hd__nor3_1 _07528_ (.A(_01405_),
    .B(_01440_),
    .C(_01441_),
    .Y(_01443_));
 sky130_fd_sc_hd__o21a_1 _07529_ (.A1(_01440_),
    .A2(_01441_),
    .B1(_01405_),
    .X(_01444_));
 sky130_fd_sc_hd__a21o_1 _07530_ (.A1(_01309_),
    .A2(_01318_),
    .B1(_01317_),
    .X(_01445_));
 sky130_fd_sc_hd__nand2_1 _07531_ (.A(net401),
    .B(net180),
    .Y(_01446_));
 sky130_fd_sc_hd__and4_1 _07532_ (.A(net414),
    .B(net406),
    .C(net173),
    .D(net165),
    .X(_01447_));
 sky130_fd_sc_hd__a22o_1 _07533_ (.A1(net406),
    .A2(net173),
    .B1(net165),
    .B2(net414),
    .X(_01448_));
 sky130_fd_sc_hd__and2b_1 _07534_ (.A_N(_01447_),
    .B(_01448_),
    .X(_01449_));
 sky130_fd_sc_hd__xnor2_1 _07535_ (.A(_01446_),
    .B(_01449_),
    .Y(_01450_));
 sky130_fd_sc_hd__and2_1 _07536_ (.A(net421),
    .B(net620),
    .X(_01451_));
 sky130_fd_sc_hd__nand4_1 _07537_ (.A(net183),
    .B(net428),
    .C(net612),
    .D(net596),
    .Y(_01452_));
 sky130_fd_sc_hd__a22o_1 _07538_ (.A1(net428),
    .A2(net612),
    .B1(net596),
    .B2(net183),
    .X(_01454_));
 sky130_fd_sc_hd__nand3_1 _07539_ (.A(_01451_),
    .B(_01452_),
    .C(_01454_),
    .Y(_01455_));
 sky130_fd_sc_hd__a21o_1 _07540_ (.A1(_01452_),
    .A2(_01454_),
    .B1(_01451_),
    .X(_01456_));
 sky130_fd_sc_hd__a31o_1 _07541_ (.A1(net421),
    .A2(net165),
    .A3(_01295_),
    .B1(_01294_),
    .X(_01457_));
 sky130_fd_sc_hd__nand3_1 _07542_ (.A(_01455_),
    .B(_01456_),
    .C(_01457_),
    .Y(_01458_));
 sky130_fd_sc_hd__a21o_1 _07543_ (.A1(_01455_),
    .A2(_01456_),
    .B1(_01457_),
    .X(_01459_));
 sky130_fd_sc_hd__nand3_1 _07544_ (.A(_01450_),
    .B(_01458_),
    .C(_01459_),
    .Y(_01460_));
 sky130_fd_sc_hd__a21o_1 _07545_ (.A1(_01458_),
    .A2(_01459_),
    .B1(_01450_),
    .X(_01461_));
 sky130_fd_sc_hd__nand3_2 _07546_ (.A(_01445_),
    .B(_01460_),
    .C(_01461_),
    .Y(_01462_));
 sky130_fd_sc_hd__a21o_1 _07547_ (.A1(_01460_),
    .A2(_01461_),
    .B1(_01445_),
    .X(_01463_));
 sky130_fd_sc_hd__o211ai_2 _07548_ (.A1(_01299_),
    .A2(_01302_),
    .B1(_01462_),
    .C1(_01463_),
    .Y(_01465_));
 sky130_fd_sc_hd__a211o_1 _07549_ (.A1(_01462_),
    .A2(_01463_),
    .B1(_01299_),
    .C1(_01302_),
    .X(_01466_));
 sky130_fd_sc_hd__nand2_1 _07550_ (.A(_01465_),
    .B(_01466_),
    .Y(_01467_));
 sky130_fd_sc_hd__nand2_1 _07551_ (.A(_01313_),
    .B(_01315_),
    .Y(_01468_));
 sky130_fd_sc_hd__o21bai_1 _07552_ (.A1(_01321_),
    .A2(_01324_),
    .B1_N(_01323_),
    .Y(_01469_));
 sky130_fd_sc_hd__nand2_1 _07553_ (.A(net193),
    .B(net589),
    .Y(_01470_));
 sky130_fd_sc_hd__nand4_1 _07554_ (.A(net209),
    .B(net202),
    .C(net581),
    .D(net575),
    .Y(_01471_));
 sky130_fd_sc_hd__a22o_1 _07555_ (.A1(net202),
    .A2(net581),
    .B1(net575),
    .B2(net209),
    .X(_01472_));
 sky130_fd_sc_hd__nand3b_1 _07556_ (.A_N(_01470_),
    .B(_01471_),
    .C(_01472_),
    .Y(_01473_));
 sky130_fd_sc_hd__a21bo_1 _07557_ (.A1(_01471_),
    .A2(_01472_),
    .B1_N(_01470_),
    .X(_01474_));
 sky130_fd_sc_hd__and3_1 _07558_ (.A(_01469_),
    .B(_01473_),
    .C(_01474_),
    .X(_01476_));
 sky130_fd_sc_hd__a21o_1 _07559_ (.A1(_01473_),
    .A2(_01474_),
    .B1(_01469_),
    .X(_01477_));
 sky130_fd_sc_hd__and2b_1 _07560_ (.A_N(_01476_),
    .B(_01477_),
    .X(_01478_));
 sky130_fd_sc_hd__xor2_2 _07561_ (.A(_01468_),
    .B(_01478_),
    .X(_01479_));
 sky130_fd_sc_hd__nand2_1 _07562_ (.A(net216),
    .B(net568),
    .Y(_01480_));
 sky130_fd_sc_hd__and4_1 _07563_ (.A(net237),
    .B(net229),
    .C(net562),
    .D(net554),
    .X(_01481_));
 sky130_fd_sc_hd__a22oi_1 _07564_ (.A1(net230),
    .A2(net562),
    .B1(net554),
    .B2(net237),
    .Y(_01482_));
 sky130_fd_sc_hd__nor2_1 _07565_ (.A(_01481_),
    .B(_01482_),
    .Y(_01483_));
 sky130_fd_sc_hd__xnor2_1 _07566_ (.A(_01480_),
    .B(_01483_),
    .Y(_01484_));
 sky130_fd_sc_hd__and2_1 _07567_ (.A(net257),
    .B(net540),
    .X(_01485_));
 sky130_fd_sc_hd__nand4_1 _07568_ (.A(net436),
    .B(net344),
    .C(net534),
    .D(net526),
    .Y(_01487_));
 sky130_fd_sc_hd__a22o_1 _07569_ (.A1(net344),
    .A2(net534),
    .B1(net526),
    .B2(net436),
    .X(_01488_));
 sky130_fd_sc_hd__nand3_1 _07570_ (.A(_01485_),
    .B(_01487_),
    .C(_01488_),
    .Y(_01489_));
 sky130_fd_sc_hd__a21o_1 _07571_ (.A1(_01487_),
    .A2(_01488_),
    .B1(_01485_),
    .X(_01490_));
 sky130_fd_sc_hd__o21bai_1 _07572_ (.A1(_01327_),
    .A2(_01329_),
    .B1_N(_01328_),
    .Y(_01491_));
 sky130_fd_sc_hd__nand3_1 _07573_ (.A(_01489_),
    .B(_01490_),
    .C(_01491_),
    .Y(_01492_));
 sky130_fd_sc_hd__a21o_1 _07574_ (.A1(_01489_),
    .A2(_01490_),
    .B1(_01491_),
    .X(_01493_));
 sky130_fd_sc_hd__nand3_1 _07575_ (.A(_01484_),
    .B(_01492_),
    .C(_01493_),
    .Y(_01494_));
 sky130_fd_sc_hd__a21o_1 _07576_ (.A1(_01492_),
    .A2(_01493_),
    .B1(_01484_),
    .X(_01495_));
 sky130_fd_sc_hd__a21bo_1 _07577_ (.A1(_01326_),
    .A2(_01335_),
    .B1_N(_01334_),
    .X(_01496_));
 sky130_fd_sc_hd__nand3_4 _07578_ (.A(_01494_),
    .B(_01495_),
    .C(_01496_),
    .Y(_01498_));
 sky130_fd_sc_hd__a21o_1 _07579_ (.A1(_01494_),
    .A2(_01495_),
    .B1(_01496_),
    .X(_01499_));
 sky130_fd_sc_hd__and3_1 _07580_ (.A(_01479_),
    .B(_01498_),
    .C(_01499_),
    .X(_01500_));
 sky130_fd_sc_hd__nand3_2 _07581_ (.A(_01479_),
    .B(_01498_),
    .C(_01499_),
    .Y(_01501_));
 sky130_fd_sc_hd__a21oi_2 _07582_ (.A1(_01498_),
    .A2(_01499_),
    .B1(_01479_),
    .Y(_01502_));
 sky130_fd_sc_hd__a211oi_4 _07583_ (.A1(_01339_),
    .A2(_01342_),
    .B1(_01500_),
    .C1(_01502_),
    .Y(_01503_));
 sky130_fd_sc_hd__o211a_1 _07584_ (.A1(_01500_),
    .A2(_01502_),
    .B1(_01339_),
    .C1(_01342_),
    .X(_01504_));
 sky130_fd_sc_hd__nor3_2 _07585_ (.A(_01467_),
    .B(_01503_),
    .C(_01504_),
    .Y(_01505_));
 sky130_fd_sc_hd__o21a_1 _07586_ (.A1(_01503_),
    .A2(_01504_),
    .B1(_01467_),
    .X(_01506_));
 sky130_fd_sc_hd__a211o_1 _07587_ (.A1(_01345_),
    .A2(_01347_),
    .B1(_01505_),
    .C1(_01506_),
    .X(_01507_));
 sky130_fd_sc_hd__o211ai_1 _07588_ (.A1(_01505_),
    .A2(_01506_),
    .B1(_01345_),
    .C1(_01347_),
    .Y(_01509_));
 sky130_fd_sc_hd__or4bb_2 _07589_ (.A(_01443_),
    .B(_01444_),
    .C_N(_01507_),
    .D_N(_01509_),
    .X(_01510_));
 sky130_fd_sc_hd__a2bb2o_1 _07590_ (.A1_N(_01443_),
    .A2_N(_01444_),
    .B1(_01507_),
    .B2(_01509_),
    .X(_01511_));
 sky130_fd_sc_hd__o211ai_2 _07591_ (.A1(_01349_),
    .A2(_01351_),
    .B1(_01510_),
    .C1(_01511_),
    .Y(_01512_));
 sky130_fd_sc_hd__a211o_1 _07592_ (.A1(_01510_),
    .A2(_01511_),
    .B1(_01349_),
    .C1(_01351_),
    .X(_01513_));
 sky130_fd_sc_hd__or4bb_2 _07593_ (.A(_01403_),
    .B(_01404_),
    .C_N(_01512_),
    .D_N(_01513_),
    .X(_01514_));
 sky130_fd_sc_hd__a2bb2o_1 _07594_ (.A1_N(_01403_),
    .A2_N(_01404_),
    .B1(_01512_),
    .B2(_01513_),
    .X(_01515_));
 sky130_fd_sc_hd__o211a_1 _07595_ (.A1(_01353_),
    .A2(_01357_),
    .B1(_01514_),
    .C1(_01515_),
    .X(_01516_));
 sky130_fd_sc_hd__a211oi_1 _07596_ (.A1(_01514_),
    .A2(_01515_),
    .B1(_01353_),
    .C1(_01357_),
    .Y(_01517_));
 sky130_fd_sc_hd__a211oi_2 _07597_ (.A1(_01245_),
    .A2(_01248_),
    .B1(_01516_),
    .C1(_01517_),
    .Y(_01518_));
 sky130_fd_sc_hd__o211a_1 _07598_ (.A1(_01516_),
    .A2(_01517_),
    .B1(_01245_),
    .C1(_01248_),
    .X(_01520_));
 sky130_fd_sc_hd__a211o_2 _07599_ (.A1(_01360_),
    .A2(_01362_),
    .B1(_01518_),
    .C1(_01520_),
    .X(_01521_));
 sky130_fd_sc_hd__o211ai_2 _07600_ (.A1(_01518_),
    .A2(_01520_),
    .B1(_01360_),
    .C1(_01362_),
    .Y(_01522_));
 sky130_fd_sc_hd__a21oi_1 _07601_ (.A1(_01521_),
    .A2(_01522_),
    .B1(_01364_),
    .Y(_01523_));
 sky130_fd_sc_hd__a21o_1 _07602_ (.A1(_01521_),
    .A2(_01522_),
    .B1(_01364_),
    .X(_01524_));
 sky130_fd_sc_hd__and3_1 _07603_ (.A(_01364_),
    .B(_01521_),
    .C(_01522_),
    .X(_01525_));
 sky130_fd_sc_hd__or2_1 _07604_ (.A(_01523_),
    .B(_01525_),
    .X(_01526_));
 sky130_fd_sc_hd__o21bai_1 _07605_ (.A1(_01217_),
    .A2(_01369_),
    .B1_N(_01367_),
    .Y(_01527_));
 sky130_fd_sc_hd__xnor2_1 _07606_ (.A(_01526_),
    .B(_01527_),
    .Y(net86));
 sky130_fd_sc_hd__nor2_1 _07607_ (.A(_01516_),
    .B(_01518_),
    .Y(_01528_));
 sky130_fd_sc_hd__and4_1 _07608_ (.A(net496),
    .B(net517),
    .C(net282),
    .D(net274),
    .X(_01530_));
 sky130_fd_sc_hd__a22oi_1 _07609_ (.A1(net497),
    .A2(net282),
    .B1(net274),
    .B2(net517),
    .Y(_01531_));
 sky130_fd_sc_hd__nor2_1 _07610_ (.A(_01530_),
    .B(_01531_),
    .Y(_01532_));
 sky130_fd_sc_hd__nand2_1 _07611_ (.A(net602),
    .B(net264),
    .Y(_01533_));
 sky130_fd_sc_hd__xnor2_1 _07612_ (.A(_01532_),
    .B(_01533_),
    .Y(_01534_));
 sky130_fd_sc_hd__o21ba_1 _07613_ (.A1(_01371_),
    .A2(_01373_),
    .B1_N(_01370_),
    .X(_01535_));
 sky130_fd_sc_hd__nand2b_1 _07614_ (.A_N(_01535_),
    .B(_01534_),
    .Y(_01536_));
 sky130_fd_sc_hd__xnor2_1 _07615_ (.A(_01534_),
    .B(_01535_),
    .Y(_01537_));
 sky130_fd_sc_hd__nand3_1 _07616_ (.A(net628),
    .B(net253),
    .C(_01537_),
    .Y(_01538_));
 sky130_fd_sc_hd__a21o_1 _07617_ (.A1(net628),
    .A2(net253),
    .B1(_01537_),
    .X(_01539_));
 sky130_fd_sc_hd__nand2_1 _07618_ (.A(_01538_),
    .B(_01539_),
    .Y(_01541_));
 sky130_fd_sc_hd__nor2_1 _07619_ (.A(_01375_),
    .B(_01541_),
    .Y(_01542_));
 sky130_fd_sc_hd__and2_1 _07620_ (.A(_01375_),
    .B(_01541_),
    .X(_01543_));
 sky130_fd_sc_hd__or2_1 _07621_ (.A(_01542_),
    .B(_01543_),
    .X(_01544_));
 sky130_fd_sc_hd__a21o_1 _07622_ (.A1(_01411_),
    .A2(_01419_),
    .B1(_01418_),
    .X(_01545_));
 sky130_fd_sc_hd__a31o_1 _07623_ (.A1(net496),
    .A2(net289),
    .A3(_01383_),
    .B1(_01381_),
    .X(_01546_));
 sky130_fd_sc_hd__a31o_1 _07624_ (.A1(net474),
    .A2(net316),
    .A3(_01407_),
    .B1(_01406_),
    .X(_01547_));
 sky130_fd_sc_hd__nand4_1 _07625_ (.A(net482),
    .B(net474),
    .C(net308),
    .D(net294),
    .Y(_01548_));
 sky130_fd_sc_hd__a22o_1 _07626_ (.A1(net474),
    .A2(net309),
    .B1(net294),
    .B2(net482),
    .X(_01549_));
 sky130_fd_sc_hd__a22o_1 _07627_ (.A1(net489),
    .A2(net289),
    .B1(_01548_),
    .B2(_01549_),
    .X(_01550_));
 sky130_fd_sc_hd__nand4_1 _07628_ (.A(net489),
    .B(net289),
    .C(_01548_),
    .D(_01549_),
    .Y(_01552_));
 sky130_fd_sc_hd__nand3_1 _07629_ (.A(_01547_),
    .B(_01550_),
    .C(_01552_),
    .Y(_01553_));
 sky130_fd_sc_hd__a21o_1 _07630_ (.A1(_01550_),
    .A2(_01552_),
    .B1(_01547_),
    .X(_01554_));
 sky130_fd_sc_hd__nand3_1 _07631_ (.A(_01546_),
    .B(_01553_),
    .C(_01554_),
    .Y(_01555_));
 sky130_fd_sc_hd__a21o_1 _07632_ (.A1(_01553_),
    .A2(_01554_),
    .B1(_01546_),
    .X(_01556_));
 sky130_fd_sc_hd__and3_1 _07633_ (.A(_01545_),
    .B(_01555_),
    .C(_01556_),
    .X(_01557_));
 sky130_fd_sc_hd__a21oi_1 _07634_ (.A1(_01555_),
    .A2(_01556_),
    .B1(_01545_),
    .Y(_01558_));
 sky130_fd_sc_hd__a211oi_2 _07635_ (.A1(_01386_),
    .A2(_01389_),
    .B1(_01557_),
    .C1(_01558_),
    .Y(_01559_));
 sky130_fd_sc_hd__inv_2 _07636_ (.A(_01559_),
    .Y(_01560_));
 sky130_fd_sc_hd__o211ai_2 _07637_ (.A1(_01557_),
    .A2(_01558_),
    .B1(_01386_),
    .C1(_01389_),
    .Y(_01561_));
 sky130_fd_sc_hd__o211a_1 _07638_ (.A1(_01391_),
    .A2(_01393_),
    .B1(_01560_),
    .C1(_01561_),
    .X(_01563_));
 sky130_fd_sc_hd__a211oi_1 _07639_ (.A1(_01560_),
    .A2(_01561_),
    .B1(_01391_),
    .C1(_01393_),
    .Y(_01564_));
 sky130_fd_sc_hd__or3_1 _07640_ (.A(_01544_),
    .B(_01563_),
    .C(_01564_),
    .X(_01565_));
 sky130_fd_sc_hd__o21ai_1 _07641_ (.A1(_01563_),
    .A2(_01564_),
    .B1(_01544_),
    .Y(_01566_));
 sky130_fd_sc_hd__o211a_1 _07642_ (.A1(_01440_),
    .A2(_01443_),
    .B1(_01565_),
    .C1(_01566_),
    .X(_01567_));
 sky130_fd_sc_hd__a211oi_1 _07643_ (.A1(_01565_),
    .A2(_01566_),
    .B1(_01440_),
    .C1(_01443_),
    .Y(_01568_));
 sky130_fd_sc_hd__a211oi_1 _07644_ (.A1(_01396_),
    .A2(_01399_),
    .B1(_01567_),
    .C1(_01568_),
    .Y(_01569_));
 sky130_fd_sc_hd__o211a_1 _07645_ (.A1(_01567_),
    .A2(_01568_),
    .B1(_01396_),
    .C1(_01399_),
    .X(_01570_));
 sky130_fd_sc_hd__and4_1 _07646_ (.A(net450),
    .B(net443),
    .C(net331),
    .D(net324),
    .X(_01571_));
 sky130_fd_sc_hd__a22o_1 _07647_ (.A1(net443),
    .A2(net331),
    .B1(net324),
    .B2(net450),
    .X(_01572_));
 sky130_fd_sc_hd__and2b_1 _07648_ (.A_N(_01571_),
    .B(_01572_),
    .X(_01574_));
 sky130_fd_sc_hd__nand2_1 _07649_ (.A(net459),
    .B(net317),
    .Y(_01575_));
 sky130_fd_sc_hd__xnor2_1 _07650_ (.A(_01574_),
    .B(_01575_),
    .Y(_01576_));
 sky130_fd_sc_hd__nand2_1 _07651_ (.A(net544),
    .B(net339),
    .Y(_01577_));
 sky130_fd_sc_hd__and4_1 _07652_ (.A(net469),
    .B(net382),
    .C(net361),
    .D(net353),
    .X(_01578_));
 sky130_fd_sc_hd__a22oi_2 _07653_ (.A1(net383),
    .A2(net361),
    .B1(net353),
    .B2(net469),
    .Y(_01579_));
 sky130_fd_sc_hd__or3_1 _07654_ (.A(_01577_),
    .B(_01578_),
    .C(_01579_),
    .X(_01580_));
 sky130_fd_sc_hd__o21ai_1 _07655_ (.A1(_01578_),
    .A2(_01579_),
    .B1(_01577_),
    .Y(_01581_));
 sky130_fd_sc_hd__o21bai_1 _07656_ (.A1(_01412_),
    .A2(_01414_),
    .B1_N(_01413_),
    .Y(_01582_));
 sky130_fd_sc_hd__and3_1 _07657_ (.A(_01580_),
    .B(_01581_),
    .C(_01582_),
    .X(_01583_));
 sky130_fd_sc_hd__a21o_1 _07658_ (.A1(_01580_),
    .A2(_01581_),
    .B1(_01582_),
    .X(_01585_));
 sky130_fd_sc_hd__and2b_1 _07659_ (.A_N(_01583_),
    .B(_01585_),
    .X(_01586_));
 sky130_fd_sc_hd__xnor2_1 _07660_ (.A(_01576_),
    .B(_01586_),
    .Y(_01587_));
 sky130_fd_sc_hd__nand2_1 _07661_ (.A(_01425_),
    .B(_01428_),
    .Y(_01588_));
 sky130_fd_sc_hd__a31o_1 _07662_ (.A1(net399),
    .A2(net180),
    .A3(_01448_),
    .B1(_01447_),
    .X(_01589_));
 sky130_fd_sc_hd__nand4_1 _07663_ (.A(net225),
    .B(net180),
    .C(net391),
    .D(net375),
    .Y(_01590_));
 sky130_fd_sc_hd__a22o_1 _07664_ (.A1(net180),
    .A2(net391),
    .B1(net375),
    .B2(net225),
    .X(_01591_));
 sky130_fd_sc_hd__a22o_1 _07665_ (.A1(net301),
    .A2(net372),
    .B1(_01590_),
    .B2(_01591_),
    .X(_01592_));
 sky130_fd_sc_hd__nand4_1 _07666_ (.A(net301),
    .B(net368),
    .C(_01590_),
    .D(_01591_),
    .Y(_01593_));
 sky130_fd_sc_hd__nand3_1 _07667_ (.A(_01589_),
    .B(_01592_),
    .C(_01593_),
    .Y(_01594_));
 sky130_fd_sc_hd__a21o_1 _07668_ (.A1(_01592_),
    .A2(_01593_),
    .B1(_01589_),
    .X(_01596_));
 sky130_fd_sc_hd__nand3_1 _07669_ (.A(_01588_),
    .B(_01594_),
    .C(_01596_),
    .Y(_01597_));
 sky130_fd_sc_hd__a21o_1 _07670_ (.A1(_01594_),
    .A2(_01596_),
    .B1(_01588_),
    .X(_01598_));
 sky130_fd_sc_hd__a21bo_1 _07671_ (.A1(_01423_),
    .A2(_01430_),
    .B1_N(_01429_),
    .X(_01599_));
 sky130_fd_sc_hd__and3_1 _07672_ (.A(_01597_),
    .B(_01598_),
    .C(_01599_),
    .X(_01600_));
 sky130_fd_sc_hd__a21oi_1 _07673_ (.A1(_01597_),
    .A2(_01598_),
    .B1(_01599_),
    .Y(_01601_));
 sky130_fd_sc_hd__nor3_1 _07674_ (.A(_01587_),
    .B(_01600_),
    .C(_01601_),
    .Y(_01602_));
 sky130_fd_sc_hd__o21a_1 _07675_ (.A1(_01600_),
    .A2(_01601_),
    .B1(_01587_),
    .X(_01603_));
 sky130_fd_sc_hd__a211oi_1 _07676_ (.A1(_01462_),
    .A2(_01465_),
    .B1(_01602_),
    .C1(_01603_),
    .Y(_01604_));
 sky130_fd_sc_hd__o211a_1 _07677_ (.A1(_01602_),
    .A2(_01603_),
    .B1(_01462_),
    .C1(_01465_),
    .X(_01605_));
 sky130_fd_sc_hd__a211oi_1 _07678_ (.A1(_01436_),
    .A2(_01438_),
    .B1(_01604_),
    .C1(_01605_),
    .Y(_01607_));
 sky130_fd_sc_hd__o211a_1 _07679_ (.A1(_01604_),
    .A2(_01605_),
    .B1(_01436_),
    .C1(_01438_),
    .X(_01608_));
 sky130_fd_sc_hd__nand2_1 _07680_ (.A(_01458_),
    .B(_01460_),
    .Y(_01609_));
 sky130_fd_sc_hd__a21o_1 _07681_ (.A1(_01468_),
    .A2(_01477_),
    .B1(_01476_),
    .X(_01610_));
 sky130_fd_sc_hd__nand2_1 _07682_ (.A(net399),
    .B(net173),
    .Y(_01611_));
 sky130_fd_sc_hd__and4_1 _07683_ (.A(net414),
    .B(net406),
    .C(net165),
    .D(net618),
    .X(_01612_));
 sky130_fd_sc_hd__a22o_1 _07684_ (.A1(net406),
    .A2(net165),
    .B1(net618),
    .B2(net414),
    .X(_01613_));
 sky130_fd_sc_hd__and2b_1 _07685_ (.A_N(_01612_),
    .B(_01613_),
    .X(_01614_));
 sky130_fd_sc_hd__xnor2_1 _07686_ (.A(_01611_),
    .B(_01614_),
    .Y(_01615_));
 sky130_fd_sc_hd__nand2_1 _07687_ (.A(net421),
    .B(net610),
    .Y(_01616_));
 sky130_fd_sc_hd__and4_1 _07688_ (.A(net182),
    .B(net428),
    .C(net594),
    .D(net587),
    .X(_01618_));
 sky130_fd_sc_hd__a22oi_2 _07689_ (.A1(net428),
    .A2(net596),
    .B1(net587),
    .B2(net183),
    .Y(_01619_));
 sky130_fd_sc_hd__or3_1 _07690_ (.A(_01616_),
    .B(_01618_),
    .C(_01619_),
    .X(_01620_));
 sky130_fd_sc_hd__o21ai_1 _07691_ (.A1(_01618_),
    .A2(_01619_),
    .B1(_01616_),
    .Y(_01621_));
 sky130_fd_sc_hd__a21bo_1 _07692_ (.A1(_01451_),
    .A2(_01454_),
    .B1_N(_01452_),
    .X(_01622_));
 sky130_fd_sc_hd__nand3_1 _07693_ (.A(_01620_),
    .B(_01621_),
    .C(_01622_),
    .Y(_01623_));
 sky130_fd_sc_hd__a21o_1 _07694_ (.A1(_01620_),
    .A2(_01621_),
    .B1(_01622_),
    .X(_01624_));
 sky130_fd_sc_hd__nand3_1 _07695_ (.A(_01615_),
    .B(_01623_),
    .C(_01624_),
    .Y(_01625_));
 sky130_fd_sc_hd__a21o_1 _07696_ (.A1(_01623_),
    .A2(_01624_),
    .B1(_01615_),
    .X(_01626_));
 sky130_fd_sc_hd__nand3_2 _07697_ (.A(_01610_),
    .B(_01625_),
    .C(_01626_),
    .Y(_01627_));
 sky130_fd_sc_hd__a21o_1 _07698_ (.A1(_01625_),
    .A2(_01626_),
    .B1(_01610_),
    .X(_01629_));
 sky130_fd_sc_hd__nand3_2 _07699_ (.A(_01609_),
    .B(_01627_),
    .C(_01629_),
    .Y(_01630_));
 sky130_fd_sc_hd__a21o_1 _07700_ (.A1(_01627_),
    .A2(_01629_),
    .B1(_01609_),
    .X(_01631_));
 sky130_fd_sc_hd__nand2_1 _07701_ (.A(_01471_),
    .B(_01473_),
    .Y(_01632_));
 sky130_fd_sc_hd__o21bai_1 _07702_ (.A1(_01480_),
    .A2(_01482_),
    .B1_N(_01481_),
    .Y(_01633_));
 sky130_fd_sc_hd__nand2_1 _07703_ (.A(net192),
    .B(net579),
    .Y(_01634_));
 sky130_fd_sc_hd__nand4_1 _07704_ (.A(net209),
    .B(net202),
    .C(net575),
    .D(net568),
    .Y(_01635_));
 sky130_fd_sc_hd__a22o_1 _07705_ (.A1(net202),
    .A2(net575),
    .B1(net568),
    .B2(net209),
    .X(_01636_));
 sky130_fd_sc_hd__nand3b_1 _07706_ (.A_N(_01634_),
    .B(_01635_),
    .C(_01636_),
    .Y(_01637_));
 sky130_fd_sc_hd__a21bo_1 _07707_ (.A1(_01635_),
    .A2(_01636_),
    .B1_N(_01634_),
    .X(_01638_));
 sky130_fd_sc_hd__and3_1 _07708_ (.A(_01633_),
    .B(_01637_),
    .C(_01638_),
    .X(_01640_));
 sky130_fd_sc_hd__a21o_1 _07709_ (.A1(_01637_),
    .A2(_01638_),
    .B1(_01633_),
    .X(_01641_));
 sky130_fd_sc_hd__and2b_1 _07710_ (.A_N(_01640_),
    .B(_01641_),
    .X(_01642_));
 sky130_fd_sc_hd__xor2_1 _07711_ (.A(_01632_),
    .B(_01642_),
    .X(_01643_));
 sky130_fd_sc_hd__nand2_1 _07712_ (.A(net216),
    .B(net562),
    .Y(_01644_));
 sky130_fd_sc_hd__and4_1 _07713_ (.A(net237),
    .B(net229),
    .C(net554),
    .D(net538),
    .X(_01645_));
 sky130_fd_sc_hd__a22oi_1 _07714_ (.A1(net230),
    .A2(net554),
    .B1(net540),
    .B2(net237),
    .Y(_01646_));
 sky130_fd_sc_hd__nor2_1 _07715_ (.A(_01645_),
    .B(_01646_),
    .Y(_01647_));
 sky130_fd_sc_hd__xnor2_1 _07716_ (.A(_01644_),
    .B(_01647_),
    .Y(_01648_));
 sky130_fd_sc_hd__nand2_1 _07717_ (.A(net257),
    .B(net534),
    .Y(_01649_));
 sky130_fd_sc_hd__nand2_1 _07718_ (.A(net343),
    .B(net509),
    .Y(_01650_));
 sky130_fd_sc_hd__and4_1 _07719_ (.A(net441),
    .B(net343),
    .C(net526),
    .D(net511),
    .X(_01651_));
 sky130_fd_sc_hd__a22oi_2 _07720_ (.A1(net343),
    .A2(net526),
    .B1(net511),
    .B2(net441),
    .Y(_01652_));
 sky130_fd_sc_hd__or3_1 _07721_ (.A(_01649_),
    .B(_01651_),
    .C(_01652_),
    .X(_01653_));
 sky130_fd_sc_hd__o21ai_1 _07722_ (.A1(_01651_),
    .A2(_01652_),
    .B1(_01649_),
    .Y(_01654_));
 sky130_fd_sc_hd__a21bo_1 _07723_ (.A1(_01485_),
    .A2(_01488_),
    .B1_N(_01487_),
    .X(_01655_));
 sky130_fd_sc_hd__nand3_1 _07724_ (.A(_01653_),
    .B(_01654_),
    .C(_01655_),
    .Y(_01656_));
 sky130_fd_sc_hd__a21o_1 _07725_ (.A1(_01653_),
    .A2(_01654_),
    .B1(_01655_),
    .X(_01657_));
 sky130_fd_sc_hd__nand3_1 _07726_ (.A(_01648_),
    .B(_01656_),
    .C(_01657_),
    .Y(_01658_));
 sky130_fd_sc_hd__a21o_1 _07727_ (.A1(_01656_),
    .A2(_01657_),
    .B1(_01648_),
    .X(_01659_));
 sky130_fd_sc_hd__a21bo_1 _07728_ (.A1(_01484_),
    .A2(_01493_),
    .B1_N(_01492_),
    .X(_01661_));
 sky130_fd_sc_hd__and3_1 _07729_ (.A(_01658_),
    .B(_01659_),
    .C(_01661_),
    .X(_01662_));
 sky130_fd_sc_hd__a21oi_1 _07730_ (.A1(_01658_),
    .A2(_01659_),
    .B1(_01661_),
    .Y(_01663_));
 sky130_fd_sc_hd__nor3b_1 _07731_ (.A(_01662_),
    .B(_01663_),
    .C_N(_01643_),
    .Y(_01664_));
 sky130_fd_sc_hd__o21ba_1 _07732_ (.A1(_01662_),
    .A2(_01663_),
    .B1_N(_01643_),
    .X(_01665_));
 sky130_fd_sc_hd__a211oi_2 _07733_ (.A1(_01498_),
    .A2(_01501_),
    .B1(net158),
    .C1(_01665_),
    .Y(_01666_));
 sky130_fd_sc_hd__a211o_1 _07734_ (.A1(_01498_),
    .A2(_01501_),
    .B1(net158),
    .C1(_01665_),
    .X(_01667_));
 sky130_fd_sc_hd__o211ai_2 _07735_ (.A1(net158),
    .A2(_01665_),
    .B1(_01498_),
    .C1(_01501_),
    .Y(_01668_));
 sky130_fd_sc_hd__and4_1 _07736_ (.A(_01630_),
    .B(_01631_),
    .C(_01667_),
    .D(_01668_),
    .X(_01669_));
 sky130_fd_sc_hd__nand4_2 _07737_ (.A(_01630_),
    .B(_01631_),
    .C(_01667_),
    .D(_01668_),
    .Y(_01670_));
 sky130_fd_sc_hd__a22o_1 _07738_ (.A1(_01630_),
    .A2(_01631_),
    .B1(_01667_),
    .B2(_01668_),
    .X(_01672_));
 sky130_fd_sc_hd__o211ai_4 _07739_ (.A1(_01503_),
    .A2(_01505_),
    .B1(_01670_),
    .C1(_01672_),
    .Y(_01673_));
 sky130_fd_sc_hd__a211o_1 _07740_ (.A1(_01670_),
    .A2(_01672_),
    .B1(_01503_),
    .C1(_01505_),
    .X(_01674_));
 sky130_fd_sc_hd__and4bb_1 _07741_ (.A_N(_01607_),
    .B_N(_01608_),
    .C(_01673_),
    .D(_01674_),
    .X(_01675_));
 sky130_fd_sc_hd__or4bb_1 _07742_ (.A(_01607_),
    .B(_01608_),
    .C_N(_01673_),
    .D_N(_01674_),
    .X(_01676_));
 sky130_fd_sc_hd__a2bb2oi_1 _07743_ (.A1_N(_01607_),
    .A2_N(_01608_),
    .B1(_01673_),
    .B2(_01674_),
    .Y(_01677_));
 sky130_fd_sc_hd__a211oi_2 _07744_ (.A1(_01507_),
    .A2(_01510_),
    .B1(_01675_),
    .C1(_01677_),
    .Y(_01678_));
 sky130_fd_sc_hd__o211a_1 _07745_ (.A1(_01675_),
    .A2(_01677_),
    .B1(_01507_),
    .C1(_01510_),
    .X(_01679_));
 sky130_fd_sc_hd__nor4_1 _07746_ (.A(_01569_),
    .B(_01570_),
    .C(_01678_),
    .D(_01679_),
    .Y(_01680_));
 sky130_fd_sc_hd__o22a_1 _07747_ (.A1(_01569_),
    .A2(_01570_),
    .B1(_01678_),
    .B2(_01679_),
    .X(_01681_));
 sky130_fd_sc_hd__a211oi_1 _07748_ (.A1(_01512_),
    .A2(_01514_),
    .B1(net132),
    .C1(_01681_),
    .Y(_01683_));
 sky130_fd_sc_hd__a211o_1 _07749_ (.A1(_01512_),
    .A2(_01514_),
    .B1(net132),
    .C1(_01681_),
    .X(_01684_));
 sky130_fd_sc_hd__o211ai_1 _07750_ (.A1(net132),
    .A2(_01681_),
    .B1(_01512_),
    .C1(_01514_),
    .Y(_01685_));
 sky130_fd_sc_hd__o211a_1 _07751_ (.A1(_01401_),
    .A2(_01403_),
    .B1(_01684_),
    .C1(_01685_),
    .X(_01686_));
 sky130_fd_sc_hd__a211oi_1 _07752_ (.A1(_01684_),
    .A2(_01685_),
    .B1(_01401_),
    .C1(_01403_),
    .Y(_01687_));
 sky130_fd_sc_hd__nor2_1 _07753_ (.A(_01686_),
    .B(_01687_),
    .Y(_01688_));
 sky130_fd_sc_hd__nand2b_1 _07754_ (.A_N(_01528_),
    .B(_01688_),
    .Y(_01689_));
 sky130_fd_sc_hd__xnor2_1 _07755_ (.A(_01528_),
    .B(_01688_),
    .Y(_01690_));
 sky130_fd_sc_hd__and2b_1 _07756_ (.A_N(_01521_),
    .B(_01690_),
    .X(_01691_));
 sky130_fd_sc_hd__xor2_2 _07757_ (.A(_01521_),
    .B(_01690_),
    .X(_01692_));
 sky130_fd_sc_hd__a21o_1 _07758_ (.A1(_01367_),
    .A2(_01524_),
    .B1(_01525_),
    .X(_01694_));
 sky130_fd_sc_hd__inv_2 _07759_ (.A(_01694_),
    .Y(_01695_));
 sky130_fd_sc_hd__or4_1 _07760_ (.A(_01367_),
    .B(_01368_),
    .C(_01523_),
    .D(_01525_),
    .X(_01696_));
 sky130_fd_sc_hd__o21a_1 _07761_ (.A1(_01217_),
    .A2(_01696_),
    .B1(_01695_),
    .X(_01697_));
 sky130_fd_sc_hd__xor2_1 _07762_ (.A(_01692_),
    .B(_01697_),
    .X(net88));
 sky130_fd_sc_hd__or2_1 _07763_ (.A(_01567_),
    .B(_01569_),
    .X(_01698_));
 sky130_fd_sc_hd__nand2b_1 _07764_ (.A_N(_01563_),
    .B(_01565_),
    .Y(_01699_));
 sky130_fd_sc_hd__or2_1 _07765_ (.A(_01604_),
    .B(_01607_),
    .X(_01700_));
 sky130_fd_sc_hd__and4_1 _07766_ (.A(net488),
    .B(net496),
    .C(net280),
    .D(net274),
    .X(_01701_));
 sky130_fd_sc_hd__a22oi_1 _07767_ (.A1(net488),
    .A2(net282),
    .B1(net274),
    .B2(net496),
    .Y(_01702_));
 sky130_fd_sc_hd__nor2_1 _07768_ (.A(_01701_),
    .B(_01702_),
    .Y(_01704_));
 sky130_fd_sc_hd__nand2_1 _07769_ (.A(net517),
    .B(net264),
    .Y(_01705_));
 sky130_fd_sc_hd__xnor2_1 _07770_ (.A(_01704_),
    .B(_01705_),
    .Y(_01706_));
 sky130_fd_sc_hd__o21ba_1 _07771_ (.A1(_01531_),
    .A2(_01533_),
    .B1_N(_01530_),
    .X(_01707_));
 sky130_fd_sc_hd__nand2b_1 _07772_ (.A_N(_01707_),
    .B(_01706_),
    .Y(_01708_));
 sky130_fd_sc_hd__xnor2_1 _07773_ (.A(_01706_),
    .B(_01707_),
    .Y(_01709_));
 sky130_fd_sc_hd__nand2_1 _07774_ (.A(net602),
    .B(net253),
    .Y(_01710_));
 sky130_fd_sc_hd__nand3_1 _07775_ (.A(net602),
    .B(net253),
    .C(_01709_),
    .Y(_01711_));
 sky130_fd_sc_hd__xor2_1 _07776_ (.A(_01709_),
    .B(_01710_),
    .X(_01712_));
 sky130_fd_sc_hd__and3_1 _07777_ (.A(_01536_),
    .B(_01538_),
    .C(_01712_),
    .X(_01713_));
 sky130_fd_sc_hd__a21oi_1 _07778_ (.A1(_01536_),
    .A2(_01538_),
    .B1(_01712_),
    .Y(_01715_));
 sky130_fd_sc_hd__nor2_1 _07779_ (.A(_01713_),
    .B(_01715_),
    .Y(_01716_));
 sky130_fd_sc_hd__nand2_1 _07780_ (.A(net628),
    .B(net248),
    .Y(_01717_));
 sky130_fd_sc_hd__xnor2_1 _07781_ (.A(_01716_),
    .B(_01717_),
    .Y(_01718_));
 sky130_fd_sc_hd__a21o_1 _07782_ (.A1(_01576_),
    .A2(_01585_),
    .B1(_01583_),
    .X(_01719_));
 sky130_fd_sc_hd__nand2_1 _07783_ (.A(_01548_),
    .B(_01552_),
    .Y(_01720_));
 sky130_fd_sc_hd__a31o_1 _07784_ (.A1(net459),
    .A2(net317),
    .A3(_01572_),
    .B1(_01571_),
    .X(_01721_));
 sky130_fd_sc_hd__nand4_1 _07785_ (.A(net473),
    .B(net458),
    .C(net309),
    .D(net295),
    .Y(_01722_));
 sky130_fd_sc_hd__a22o_1 _07786_ (.A1(net458),
    .A2(net309),
    .B1(net295),
    .B2(net473),
    .X(_01723_));
 sky130_fd_sc_hd__a22o_1 _07787_ (.A1(net481),
    .A2(net287),
    .B1(_01722_),
    .B2(_01723_),
    .X(_01724_));
 sky130_fd_sc_hd__nand4_1 _07788_ (.A(net481),
    .B(net287),
    .C(_01722_),
    .D(_01723_),
    .Y(_01726_));
 sky130_fd_sc_hd__nand3_1 _07789_ (.A(_01721_),
    .B(_01724_),
    .C(_01726_),
    .Y(_01727_));
 sky130_fd_sc_hd__a21o_1 _07790_ (.A1(_01724_),
    .A2(_01726_),
    .B1(_01721_),
    .X(_01728_));
 sky130_fd_sc_hd__nand3_1 _07791_ (.A(_01720_),
    .B(_01727_),
    .C(_01728_),
    .Y(_01729_));
 sky130_fd_sc_hd__a21o_1 _07792_ (.A1(_01727_),
    .A2(_01728_),
    .B1(_01720_),
    .X(_01730_));
 sky130_fd_sc_hd__and3_1 _07793_ (.A(_01719_),
    .B(_01729_),
    .C(_01730_),
    .X(_01731_));
 sky130_fd_sc_hd__a21oi_1 _07794_ (.A1(_01729_),
    .A2(_01730_),
    .B1(_01719_),
    .Y(_01732_));
 sky130_fd_sc_hd__a211oi_1 _07795_ (.A1(_01553_),
    .A2(_01555_),
    .B1(_01731_),
    .C1(_01732_),
    .Y(_01733_));
 sky130_fd_sc_hd__o211a_1 _07796_ (.A1(_01731_),
    .A2(_01732_),
    .B1(_01553_),
    .C1(_01555_),
    .X(_01734_));
 sky130_fd_sc_hd__or2_1 _07797_ (.A(_01733_),
    .B(_01734_),
    .X(_01735_));
 sky130_fd_sc_hd__nor2_1 _07798_ (.A(_01557_),
    .B(_01559_),
    .Y(_01737_));
 sky130_fd_sc_hd__or2_1 _07799_ (.A(_01735_),
    .B(_01737_),
    .X(_01738_));
 sky130_fd_sc_hd__nand2_1 _07800_ (.A(_01735_),
    .B(_01737_),
    .Y(_01739_));
 sky130_fd_sc_hd__xnor2_1 _07801_ (.A(_01735_),
    .B(_01737_),
    .Y(_01740_));
 sky130_fd_sc_hd__xnor2_1 _07802_ (.A(_01718_),
    .B(_01740_),
    .Y(_01741_));
 sky130_fd_sc_hd__nand2_1 _07803_ (.A(_01700_),
    .B(_01741_),
    .Y(_01742_));
 sky130_fd_sc_hd__xor2_1 _07804_ (.A(_01700_),
    .B(_01741_),
    .X(_01743_));
 sky130_fd_sc_hd__xor2_1 _07805_ (.A(_01699_),
    .B(_01743_),
    .X(_01744_));
 sky130_fd_sc_hd__nor2_1 _07806_ (.A(_01600_),
    .B(_01602_),
    .Y(_01745_));
 sky130_fd_sc_hd__and4_1 _07807_ (.A(net544),
    .B(net443),
    .C(net331),
    .D(net324),
    .X(_01746_));
 sky130_fd_sc_hd__a22o_1 _07808_ (.A1(net544),
    .A2(net331),
    .B1(net324),
    .B2(net443),
    .X(_01748_));
 sky130_fd_sc_hd__and2b_1 _07809_ (.A_N(_01746_),
    .B(_01748_),
    .X(_01749_));
 sky130_fd_sc_hd__nand2_1 _07810_ (.A(net450),
    .B(net317),
    .Y(_01750_));
 sky130_fd_sc_hd__xnor2_1 _07811_ (.A(_01749_),
    .B(_01750_),
    .Y(_01751_));
 sky130_fd_sc_hd__nand2_1 _07812_ (.A(net469),
    .B(net339),
    .Y(_01752_));
 sky130_fd_sc_hd__and4_1 _07813_ (.A(net383),
    .B(net298),
    .C(net361),
    .D(net353),
    .X(_01753_));
 sky130_fd_sc_hd__a22oi_2 _07814_ (.A1(net298),
    .A2(net361),
    .B1(net353),
    .B2(net383),
    .Y(_01754_));
 sky130_fd_sc_hd__or3_1 _07815_ (.A(_01752_),
    .B(_01753_),
    .C(_01754_),
    .X(_01755_));
 sky130_fd_sc_hd__o21ai_1 _07816_ (.A1(_01753_),
    .A2(_01754_),
    .B1(_01752_),
    .Y(_01756_));
 sky130_fd_sc_hd__o21bai_1 _07817_ (.A1(_01577_),
    .A2(_01579_),
    .B1_N(_01578_),
    .Y(_01757_));
 sky130_fd_sc_hd__and3_1 _07818_ (.A(_01755_),
    .B(_01756_),
    .C(_01757_),
    .X(_01759_));
 sky130_fd_sc_hd__a21o_1 _07819_ (.A1(_01755_),
    .A2(_01756_),
    .B1(_01757_),
    .X(_01760_));
 sky130_fd_sc_hd__and2b_1 _07820_ (.A_N(_01759_),
    .B(_01760_),
    .X(_01761_));
 sky130_fd_sc_hd__xnor2_1 _07821_ (.A(_01751_),
    .B(_01761_),
    .Y(_01762_));
 sky130_fd_sc_hd__nand2_1 _07822_ (.A(_01590_),
    .B(_01593_),
    .Y(_01763_));
 sky130_fd_sc_hd__a31o_1 _07823_ (.A1(net399),
    .A2(net173),
    .A3(_01613_),
    .B1(_01612_),
    .X(_01764_));
 sky130_fd_sc_hd__nand4_1 _07824_ (.A(net177),
    .B(net391),
    .C(net169),
    .D(net375),
    .Y(_01765_));
 sky130_fd_sc_hd__a22o_1 _07825_ (.A1(net391),
    .A2(net169),
    .B1(net375),
    .B2(net178),
    .X(_01766_));
 sky130_fd_sc_hd__a22o_1 _07826_ (.A1(net222),
    .A2(net368),
    .B1(_01765_),
    .B2(_01766_),
    .X(_01767_));
 sky130_fd_sc_hd__nand4_1 _07827_ (.A(net222),
    .B(net368),
    .C(_01765_),
    .D(_01766_),
    .Y(_01768_));
 sky130_fd_sc_hd__nand3_1 _07828_ (.A(_01764_),
    .B(_01767_),
    .C(_01768_),
    .Y(_01770_));
 sky130_fd_sc_hd__a21o_1 _07829_ (.A1(_01767_),
    .A2(_01768_),
    .B1(_01764_),
    .X(_01771_));
 sky130_fd_sc_hd__nand3_1 _07830_ (.A(_01763_),
    .B(_01770_),
    .C(_01771_),
    .Y(_01772_));
 sky130_fd_sc_hd__a21o_1 _07831_ (.A1(_01770_),
    .A2(_01771_),
    .B1(_01763_),
    .X(_01773_));
 sky130_fd_sc_hd__a21bo_1 _07832_ (.A1(_01588_),
    .A2(_01596_),
    .B1_N(_01594_),
    .X(_01774_));
 sky130_fd_sc_hd__and3_1 _07833_ (.A(_01772_),
    .B(_01773_),
    .C(_01774_),
    .X(_01775_));
 sky130_fd_sc_hd__a21oi_1 _07834_ (.A1(_01772_),
    .A2(_01773_),
    .B1(_01774_),
    .Y(_01776_));
 sky130_fd_sc_hd__nor3_1 _07835_ (.A(_01762_),
    .B(_01775_),
    .C(_01776_),
    .Y(_01777_));
 sky130_fd_sc_hd__o21a_1 _07836_ (.A1(_01775_),
    .A2(_01776_),
    .B1(_01762_),
    .X(_01778_));
 sky130_fd_sc_hd__a211oi_1 _07837_ (.A1(_01627_),
    .A2(_01630_),
    .B1(_01777_),
    .C1(_01778_),
    .Y(_01779_));
 sky130_fd_sc_hd__o211a_1 _07838_ (.A1(_01777_),
    .A2(_01778_),
    .B1(_01627_),
    .C1(_01630_),
    .X(_01781_));
 sky130_fd_sc_hd__nor2_1 _07839_ (.A(_01779_),
    .B(_01781_),
    .Y(_01782_));
 sky130_fd_sc_hd__xnor2_1 _07840_ (.A(_01745_),
    .B(_01782_),
    .Y(_01783_));
 sky130_fd_sc_hd__nand2_1 _07841_ (.A(_01623_),
    .B(_01625_),
    .Y(_01784_));
 sky130_fd_sc_hd__a21o_1 _07842_ (.A1(_01632_),
    .A2(_01641_),
    .B1(_01640_),
    .X(_01785_));
 sky130_fd_sc_hd__nand2_1 _07843_ (.A(net399),
    .B(net161),
    .Y(_01786_));
 sky130_fd_sc_hd__and4_1 _07844_ (.A(net415),
    .B(net407),
    .C(net618),
    .D(net610),
    .X(_01787_));
 sky130_fd_sc_hd__a22o_1 _07845_ (.A1(net407),
    .A2(net618),
    .B1(net610),
    .B2(net415),
    .X(_01788_));
 sky130_fd_sc_hd__and2b_1 _07846_ (.A_N(_01787_),
    .B(_01788_),
    .X(_01789_));
 sky130_fd_sc_hd__xnor2_1 _07847_ (.A(_01786_),
    .B(_01789_),
    .Y(_01790_));
 sky130_fd_sc_hd__nand2_1 _07848_ (.A(net421),
    .B(net594),
    .Y(_01792_));
 sky130_fd_sc_hd__and4_1 _07849_ (.A(net182),
    .B(net427),
    .C(net588),
    .D(net579),
    .X(_01793_));
 sky130_fd_sc_hd__a22oi_2 _07850_ (.A1(net427),
    .A2(net588),
    .B1(net579),
    .B2(net182),
    .Y(_01794_));
 sky130_fd_sc_hd__or3_1 _07851_ (.A(_01792_),
    .B(_01793_),
    .C(_01794_),
    .X(_01795_));
 sky130_fd_sc_hd__o21ai_1 _07852_ (.A1(_01793_),
    .A2(_01794_),
    .B1(_01792_),
    .Y(_01796_));
 sky130_fd_sc_hd__o21bai_1 _07853_ (.A1(_01616_),
    .A2(_01619_),
    .B1_N(_01618_),
    .Y(_01797_));
 sky130_fd_sc_hd__nand3_1 _07854_ (.A(_01795_),
    .B(_01796_),
    .C(_01797_),
    .Y(_01798_));
 sky130_fd_sc_hd__a21o_1 _07855_ (.A1(_01795_),
    .A2(_01796_),
    .B1(_01797_),
    .X(_01799_));
 sky130_fd_sc_hd__nand3_1 _07856_ (.A(_01790_),
    .B(_01798_),
    .C(_01799_),
    .Y(_01800_));
 sky130_fd_sc_hd__a21o_1 _07857_ (.A1(_01798_),
    .A2(_01799_),
    .B1(_01790_),
    .X(_01801_));
 sky130_fd_sc_hd__nand3_1 _07858_ (.A(_01785_),
    .B(_01800_),
    .C(_01801_),
    .Y(_01803_));
 sky130_fd_sc_hd__a21o_1 _07859_ (.A1(_01800_),
    .A2(_01801_),
    .B1(_01785_),
    .X(_01804_));
 sky130_fd_sc_hd__nand3_1 _07860_ (.A(_01784_),
    .B(_01803_),
    .C(_01804_),
    .Y(_01805_));
 sky130_fd_sc_hd__a21o_1 _07861_ (.A1(_01803_),
    .A2(_01804_),
    .B1(_01784_),
    .X(_01806_));
 sky130_fd_sc_hd__and2_1 _07862_ (.A(_01805_),
    .B(_01806_),
    .X(_01807_));
 sky130_fd_sc_hd__nand2_1 _07863_ (.A(_01635_),
    .B(_01637_),
    .Y(_01808_));
 sky130_fd_sc_hd__o21bai_1 _07864_ (.A1(_01644_),
    .A2(_01646_),
    .B1_N(_01645_),
    .Y(_01809_));
 sky130_fd_sc_hd__a22o_1 _07865_ (.A1(net201),
    .A2(net566),
    .B1(net559),
    .B2(net209),
    .X(_01810_));
 sky130_fd_sc_hd__nand4_1 _07866_ (.A(net209),
    .B(net201),
    .C(net566),
    .D(net559),
    .Y(_01811_));
 sky130_fd_sc_hd__a22o_1 _07867_ (.A1(net192),
    .A2(net573),
    .B1(_01810_),
    .B2(_01811_),
    .X(_01812_));
 sky130_fd_sc_hd__nand4_1 _07868_ (.A(net192),
    .B(net573),
    .C(_01810_),
    .D(_01811_),
    .Y(_01814_));
 sky130_fd_sc_hd__and3_1 _07869_ (.A(_01809_),
    .B(_01812_),
    .C(_01814_),
    .X(_01815_));
 sky130_fd_sc_hd__a21o_1 _07870_ (.A1(_01812_),
    .A2(_01814_),
    .B1(_01809_),
    .X(_01816_));
 sky130_fd_sc_hd__and2b_1 _07871_ (.A_N(_01815_),
    .B(_01816_),
    .X(_01817_));
 sky130_fd_sc_hd__xor2_1 _07872_ (.A(_01808_),
    .B(_01817_),
    .X(_01818_));
 sky130_fd_sc_hd__nand2_1 _07873_ (.A(net216),
    .B(net552),
    .Y(_01819_));
 sky130_fd_sc_hd__and4_1 _07874_ (.A(net237),
    .B(net229),
    .C(net538),
    .D(net532),
    .X(_01820_));
 sky130_fd_sc_hd__a22oi_1 _07875_ (.A1(net229),
    .A2(net538),
    .B1(net532),
    .B2(net237),
    .Y(_01821_));
 sky130_fd_sc_hd__nor2_1 _07876_ (.A(_01820_),
    .B(_01821_),
    .Y(_01822_));
 sky130_fd_sc_hd__xnor2_1 _07877_ (.A(_01819_),
    .B(_01822_),
    .Y(_01823_));
 sky130_fd_sc_hd__and2_1 _07878_ (.A(net257),
    .B(net526),
    .X(_01825_));
 sky130_fd_sc_hd__a22o_1 _07879_ (.A1(net343),
    .A2(net511),
    .B1(net504),
    .B2(net436),
    .X(_01826_));
 sky130_fd_sc_hd__nand4_1 _07880_ (.A(net436),
    .B(net343),
    .C(net512),
    .D(net504),
    .Y(_01827_));
 sky130_fd_sc_hd__nand3_1 _07881_ (.A(_01825_),
    .B(_01826_),
    .C(_01827_),
    .Y(_01828_));
 sky130_fd_sc_hd__a21o_1 _07882_ (.A1(_01826_),
    .A2(_01827_),
    .B1(_01825_),
    .X(_01829_));
 sky130_fd_sc_hd__o21bai_1 _07883_ (.A1(_01649_),
    .A2(_01652_),
    .B1_N(_01651_),
    .Y(_01830_));
 sky130_fd_sc_hd__nand3_1 _07884_ (.A(_01828_),
    .B(_01829_),
    .C(_01830_),
    .Y(_01831_));
 sky130_fd_sc_hd__a21o_1 _07885_ (.A1(_01828_),
    .A2(_01829_),
    .B1(_01830_),
    .X(_01832_));
 sky130_fd_sc_hd__nand3_1 _07886_ (.A(_01823_),
    .B(_01831_),
    .C(_01832_),
    .Y(_01833_));
 sky130_fd_sc_hd__a21o_1 _07887_ (.A1(_01831_),
    .A2(_01832_),
    .B1(_01823_),
    .X(_01834_));
 sky130_fd_sc_hd__a21bo_1 _07888_ (.A1(_01648_),
    .A2(_01657_),
    .B1_N(_01656_),
    .X(_01836_));
 sky130_fd_sc_hd__nand3_1 _07889_ (.A(_01833_),
    .B(_01834_),
    .C(_01836_),
    .Y(_01837_));
 sky130_fd_sc_hd__a21o_1 _07890_ (.A1(_01833_),
    .A2(_01834_),
    .B1(_01836_),
    .X(_01838_));
 sky130_fd_sc_hd__nand3_1 _07891_ (.A(_01818_),
    .B(_01837_),
    .C(_01838_),
    .Y(_01839_));
 sky130_fd_sc_hd__a21o_1 _07892_ (.A1(_01837_),
    .A2(_01838_),
    .B1(_01818_),
    .X(_01840_));
 sky130_fd_sc_hd__o211ai_2 _07893_ (.A1(_01662_),
    .A2(_01664_),
    .B1(_01839_),
    .C1(_01840_),
    .Y(_01841_));
 sky130_fd_sc_hd__a211o_1 _07894_ (.A1(_01839_),
    .A2(_01840_),
    .B1(_01662_),
    .C1(_01664_),
    .X(_01842_));
 sky130_fd_sc_hd__nand3_1 _07895_ (.A(_01807_),
    .B(_01841_),
    .C(_01842_),
    .Y(_01843_));
 sky130_fd_sc_hd__a21o_1 _07896_ (.A1(_01841_),
    .A2(_01842_),
    .B1(_01807_),
    .X(_01844_));
 sky130_fd_sc_hd__o211ai_2 _07897_ (.A1(_01666_),
    .A2(_01669_),
    .B1(_01843_),
    .C1(_01844_),
    .Y(_01845_));
 sky130_fd_sc_hd__a211o_1 _07898_ (.A1(_01843_),
    .A2(_01844_),
    .B1(_01666_),
    .C1(_01669_),
    .X(_01847_));
 sky130_fd_sc_hd__and3_1 _07899_ (.A(_01783_),
    .B(_01845_),
    .C(_01847_),
    .X(_01848_));
 sky130_fd_sc_hd__a21oi_1 _07900_ (.A1(_01845_),
    .A2(_01847_),
    .B1(_01783_),
    .Y(_01849_));
 sky130_fd_sc_hd__a211o_1 _07901_ (.A1(_01673_),
    .A2(_01676_),
    .B1(_01848_),
    .C1(_01849_),
    .X(_01850_));
 sky130_fd_sc_hd__o211ai_2 _07902_ (.A1(_01848_),
    .A2(_01849_),
    .B1(_01673_),
    .C1(_01676_),
    .Y(_01851_));
 sky130_fd_sc_hd__nand3_1 _07903_ (.A(_01744_),
    .B(_01850_),
    .C(_01851_),
    .Y(_01852_));
 sky130_fd_sc_hd__a21o_1 _07904_ (.A1(_01850_),
    .A2(_01851_),
    .B1(_01744_),
    .X(_01853_));
 sky130_fd_sc_hd__o211ai_2 _07905_ (.A1(_01678_),
    .A2(_01680_),
    .B1(_01852_),
    .C1(_01853_),
    .Y(_01854_));
 sky130_fd_sc_hd__a211o_1 _07906_ (.A1(_01852_),
    .A2(_01853_),
    .B1(_01678_),
    .C1(_01680_),
    .X(_01855_));
 sky130_fd_sc_hd__nand3_1 _07907_ (.A(_01698_),
    .B(_01854_),
    .C(_01855_),
    .Y(_01856_));
 sky130_fd_sc_hd__a21o_1 _07908_ (.A1(_01854_),
    .A2(_01855_),
    .B1(_01698_),
    .X(_01858_));
 sky130_fd_sc_hd__o211ai_1 _07909_ (.A1(_01683_),
    .A2(_01686_),
    .B1(_01856_),
    .C1(_01858_),
    .Y(_01859_));
 sky130_fd_sc_hd__a211o_1 _07910_ (.A1(_01856_),
    .A2(_01858_),
    .B1(_01683_),
    .C1(_01686_),
    .X(_01860_));
 sky130_fd_sc_hd__and3_1 _07911_ (.A(_01542_),
    .B(_01859_),
    .C(_01860_),
    .X(_01861_));
 sky130_fd_sc_hd__a21oi_1 _07912_ (.A1(_01859_),
    .A2(_01860_),
    .B1(_01542_),
    .Y(_01862_));
 sky130_fd_sc_hd__o21ai_1 _07913_ (.A1(_01861_),
    .A2(_01862_),
    .B1(_01689_),
    .Y(_01863_));
 sky130_fd_sc_hd__or3_1 _07914_ (.A(_01689_),
    .B(_01861_),
    .C(_01862_),
    .X(_01864_));
 sky130_fd_sc_hd__nand2_1 _07915_ (.A(_01863_),
    .B(_01864_),
    .Y(_01865_));
 sky130_fd_sc_hd__o21bai_1 _07916_ (.A1(_01692_),
    .A2(_01697_),
    .B1_N(_01691_),
    .Y(_01866_));
 sky130_fd_sc_hd__xnor2_1 _07917_ (.A(_01865_),
    .B(_01866_),
    .Y(net89));
 sky130_fd_sc_hd__a31o_1 _07918_ (.A1(net628),
    .A2(net248),
    .A3(_01716_),
    .B1(_01715_),
    .X(_01868_));
 sky130_fd_sc_hd__a21bo_1 _07919_ (.A1(_01699_),
    .A2(_01743_),
    .B1_N(_01742_),
    .X(_01869_));
 sky130_fd_sc_hd__inv_2 _07920_ (.A(_01869_),
    .Y(_01870_));
 sky130_fd_sc_hd__a21bo_1 _07921_ (.A1(_01718_),
    .A2(_01739_),
    .B1_N(_01738_),
    .X(_01871_));
 sky130_fd_sc_hd__o21bai_1 _07922_ (.A1(_01745_),
    .A2(_01781_),
    .B1_N(_01779_),
    .Y(_01872_));
 sky130_fd_sc_hd__and4_1 _07923_ (.A(net481),
    .B(net488),
    .C(net280),
    .D(net272),
    .X(_01873_));
 sky130_fd_sc_hd__a22oi_1 _07924_ (.A1(net482),
    .A2(net280),
    .B1(net272),
    .B2(net488),
    .Y(_01874_));
 sky130_fd_sc_hd__nor2_1 _07925_ (.A(_01873_),
    .B(_01874_),
    .Y(_01875_));
 sky130_fd_sc_hd__nand2_1 _07926_ (.A(net496),
    .B(net263),
    .Y(_01876_));
 sky130_fd_sc_hd__xnor2_1 _07927_ (.A(_01875_),
    .B(_01876_),
    .Y(_01877_));
 sky130_fd_sc_hd__o21ba_1 _07928_ (.A1(_01702_),
    .A2(_01705_),
    .B1_N(_01701_),
    .X(_01879_));
 sky130_fd_sc_hd__nand2b_1 _07929_ (.A_N(_01879_),
    .B(_01877_),
    .Y(_01880_));
 sky130_fd_sc_hd__xnor2_1 _07930_ (.A(_01877_),
    .B(_01879_),
    .Y(_01881_));
 sky130_fd_sc_hd__nand2_1 _07931_ (.A(net517),
    .B(net253),
    .Y(_01882_));
 sky130_fd_sc_hd__nand3_1 _07932_ (.A(net517),
    .B(net253),
    .C(_01881_),
    .Y(_01883_));
 sky130_fd_sc_hd__xor2_1 _07933_ (.A(_01881_),
    .B(_01882_),
    .X(_01884_));
 sky130_fd_sc_hd__and3_1 _07934_ (.A(_01708_),
    .B(_01711_),
    .C(_01884_),
    .X(_01885_));
 sky130_fd_sc_hd__a21oi_1 _07935_ (.A1(_01708_),
    .A2(_01711_),
    .B1(_01884_),
    .Y(_01886_));
 sky130_fd_sc_hd__nor2_1 _07936_ (.A(_01885_),
    .B(_01886_),
    .Y(_01887_));
 sky130_fd_sc_hd__nand2_1 _07937_ (.A(net602),
    .B(net248),
    .Y(_01888_));
 sky130_fd_sc_hd__xnor2_1 _07938_ (.A(_01887_),
    .B(_01888_),
    .Y(_01890_));
 sky130_fd_sc_hd__a21o_1 _07939_ (.A1(_01751_),
    .A2(_01760_),
    .B1(_01759_),
    .X(_01891_));
 sky130_fd_sc_hd__nand2_1 _07940_ (.A(_01722_),
    .B(_01726_),
    .Y(_01892_));
 sky130_fd_sc_hd__a31o_1 _07941_ (.A1(net449),
    .A2(net317),
    .A3(_01748_),
    .B1(_01746_),
    .X(_01893_));
 sky130_fd_sc_hd__nand4_1 _07942_ (.A(net458),
    .B(net449),
    .C(net309),
    .D(net295),
    .Y(_01894_));
 sky130_fd_sc_hd__a22o_1 _07943_ (.A1(net449),
    .A2(net309),
    .B1(net295),
    .B2(net458),
    .X(_01895_));
 sky130_fd_sc_hd__a22o_1 _07944_ (.A1(net473),
    .A2(net288),
    .B1(_01894_),
    .B2(_01895_),
    .X(_01896_));
 sky130_fd_sc_hd__nand4_1 _07945_ (.A(net474),
    .B(net288),
    .C(_01894_),
    .D(_01895_),
    .Y(_01897_));
 sky130_fd_sc_hd__nand3_1 _07946_ (.A(_01893_),
    .B(_01896_),
    .C(_01897_),
    .Y(_01898_));
 sky130_fd_sc_hd__a21o_1 _07947_ (.A1(_01896_),
    .A2(_01897_),
    .B1(_01893_),
    .X(_01899_));
 sky130_fd_sc_hd__nand3_1 _07948_ (.A(_01892_),
    .B(_01898_),
    .C(_01899_),
    .Y(_01901_));
 sky130_fd_sc_hd__a21o_1 _07949_ (.A1(_01898_),
    .A2(_01899_),
    .B1(_01892_),
    .X(_01902_));
 sky130_fd_sc_hd__and3_1 _07950_ (.A(_01891_),
    .B(_01901_),
    .C(_01902_),
    .X(_01903_));
 sky130_fd_sc_hd__a21oi_1 _07951_ (.A1(_01901_),
    .A2(_01902_),
    .B1(_01891_),
    .Y(_01904_));
 sky130_fd_sc_hd__a211oi_1 _07952_ (.A1(_01727_),
    .A2(_01729_),
    .B1(_01903_),
    .C1(_01904_),
    .Y(_01905_));
 sky130_fd_sc_hd__o211a_1 _07953_ (.A1(_01903_),
    .A2(_01904_),
    .B1(_01727_),
    .C1(_01729_),
    .X(_01906_));
 sky130_fd_sc_hd__or2_1 _07954_ (.A(_01905_),
    .B(_01906_),
    .X(_01907_));
 sky130_fd_sc_hd__nor2_1 _07955_ (.A(_01731_),
    .B(_01733_),
    .Y(_01908_));
 sky130_fd_sc_hd__or2_1 _07956_ (.A(_01907_),
    .B(_01908_),
    .X(_01909_));
 sky130_fd_sc_hd__nand2_1 _07957_ (.A(_01907_),
    .B(_01908_),
    .Y(_01910_));
 sky130_fd_sc_hd__xnor2_1 _07958_ (.A(_01907_),
    .B(_01908_),
    .Y(_01912_));
 sky130_fd_sc_hd__xor2_1 _07959_ (.A(_01890_),
    .B(_01912_),
    .X(_01913_));
 sky130_fd_sc_hd__nand2b_1 _07960_ (.A_N(_01913_),
    .B(_01872_),
    .Y(_01914_));
 sky130_fd_sc_hd__xor2_1 _07961_ (.A(_01872_),
    .B(_01913_),
    .X(_01915_));
 sky130_fd_sc_hd__nand2b_1 _07962_ (.A_N(_01915_),
    .B(_01871_),
    .Y(_01916_));
 sky130_fd_sc_hd__xnor2_1 _07963_ (.A(_01871_),
    .B(_01915_),
    .Y(_01917_));
 sky130_fd_sc_hd__nor2_1 _07964_ (.A(_01775_),
    .B(_01777_),
    .Y(_01918_));
 sky130_fd_sc_hd__and4_1 _07965_ (.A(net544),
    .B(net463),
    .C(net331),
    .D(net324),
    .X(_01919_));
 sky130_fd_sc_hd__a22o_1 _07966_ (.A1(net463),
    .A2(net331),
    .B1(net324),
    .B2(net544),
    .X(_01920_));
 sky130_fd_sc_hd__and2b_1 _07967_ (.A_N(_01919_),
    .B(_01920_),
    .X(_01921_));
 sky130_fd_sc_hd__nand2_1 _07968_ (.A(net442),
    .B(net317),
    .Y(_01923_));
 sky130_fd_sc_hd__xnor2_1 _07969_ (.A(_01921_),
    .B(_01923_),
    .Y(_01924_));
 sky130_fd_sc_hd__nand4_1 _07970_ (.A(net299),
    .B(net222),
    .C(net361),
    .D(net353),
    .Y(_01925_));
 sky130_fd_sc_hd__a22o_1 _07971_ (.A1(net222),
    .A2(net361),
    .B1(net353),
    .B2(net299),
    .X(_01926_));
 sky130_fd_sc_hd__and2_1 _07972_ (.A(net383),
    .B(net339),
    .X(_01927_));
 sky130_fd_sc_hd__a21o_1 _07973_ (.A1(_01925_),
    .A2(_01926_),
    .B1(_01927_),
    .X(_01928_));
 sky130_fd_sc_hd__nand3_1 _07974_ (.A(_01925_),
    .B(_01926_),
    .C(_01927_),
    .Y(_01929_));
 sky130_fd_sc_hd__o21bai_1 _07975_ (.A1(_01752_),
    .A2(_01754_),
    .B1_N(_01753_),
    .Y(_01930_));
 sky130_fd_sc_hd__and3_1 _07976_ (.A(_01928_),
    .B(_01929_),
    .C(_01930_),
    .X(_01931_));
 sky130_fd_sc_hd__a21o_1 _07977_ (.A1(_01928_),
    .A2(_01929_),
    .B1(_01930_),
    .X(_01932_));
 sky130_fd_sc_hd__and2b_1 _07978_ (.A_N(_01931_),
    .B(_01932_),
    .X(_01934_));
 sky130_fd_sc_hd__xnor2_1 _07979_ (.A(_01924_),
    .B(_01934_),
    .Y(_01935_));
 sky130_fd_sc_hd__nand2_1 _07980_ (.A(_01765_),
    .B(_01768_),
    .Y(_01936_));
 sky130_fd_sc_hd__a31o_1 _07981_ (.A1(net400),
    .A2(net161),
    .A3(_01788_),
    .B1(_01787_),
    .X(_01937_));
 sky130_fd_sc_hd__nand4_1 _07982_ (.A(net391),
    .B(net169),
    .C(net375),
    .D(net161),
    .Y(_01938_));
 sky130_fd_sc_hd__a22o_1 _07983_ (.A1(net170),
    .A2(net376),
    .B1(net162),
    .B2(net392),
    .X(_01939_));
 sky130_fd_sc_hd__a22o_1 _07984_ (.A1(net178),
    .A2(net368),
    .B1(_01938_),
    .B2(_01939_),
    .X(_01940_));
 sky130_fd_sc_hd__nand4_1 _07985_ (.A(net178),
    .B(net368),
    .C(_01938_),
    .D(_01939_),
    .Y(_01941_));
 sky130_fd_sc_hd__nand3_1 _07986_ (.A(_01937_),
    .B(_01940_),
    .C(_01941_),
    .Y(_01942_));
 sky130_fd_sc_hd__a21o_1 _07987_ (.A1(_01940_),
    .A2(_01941_),
    .B1(_01937_),
    .X(_01943_));
 sky130_fd_sc_hd__nand3_1 _07988_ (.A(_01936_),
    .B(_01942_),
    .C(_01943_),
    .Y(_01945_));
 sky130_fd_sc_hd__a21o_1 _07989_ (.A1(_01942_),
    .A2(_01943_),
    .B1(_01936_),
    .X(_01946_));
 sky130_fd_sc_hd__a21bo_1 _07990_ (.A1(_01763_),
    .A2(_01771_),
    .B1_N(_01770_),
    .X(_01947_));
 sky130_fd_sc_hd__and3_1 _07991_ (.A(_01945_),
    .B(_01946_),
    .C(_01947_),
    .X(_01948_));
 sky130_fd_sc_hd__a21oi_1 _07992_ (.A1(_01945_),
    .A2(_01946_),
    .B1(_01947_),
    .Y(_01949_));
 sky130_fd_sc_hd__nor3_1 _07993_ (.A(_01935_),
    .B(_01948_),
    .C(_01949_),
    .Y(_01950_));
 sky130_fd_sc_hd__o21a_1 _07994_ (.A1(_01948_),
    .A2(_01949_),
    .B1(_01935_),
    .X(_01951_));
 sky130_fd_sc_hd__a211o_1 _07995_ (.A1(_01803_),
    .A2(_01805_),
    .B1(_01950_),
    .C1(_01951_),
    .X(_01952_));
 sky130_fd_sc_hd__o211ai_1 _07996_ (.A1(_01950_),
    .A2(_01951_),
    .B1(_01803_),
    .C1(_01805_),
    .Y(_01953_));
 sky130_fd_sc_hd__nand2_1 _07997_ (.A(_01952_),
    .B(_01953_),
    .Y(_01954_));
 sky130_fd_sc_hd__xor2_1 _07998_ (.A(_01918_),
    .B(_01954_),
    .X(_01956_));
 sky130_fd_sc_hd__a21o_1 _07999_ (.A1(_01808_),
    .A2(_01816_),
    .B1(_01815_),
    .X(_01957_));
 sky130_fd_sc_hd__and4_1 _08000_ (.A(net415),
    .B(net407),
    .C(net610),
    .D(net594),
    .X(_01958_));
 sky130_fd_sc_hd__a22o_1 _08001_ (.A1(net407),
    .A2(net610),
    .B1(net594),
    .B2(net415),
    .X(_01959_));
 sky130_fd_sc_hd__and2b_1 _08002_ (.A_N(_01958_),
    .B(_01959_),
    .X(_01960_));
 sky130_fd_sc_hd__nand2_1 _08003_ (.A(net400),
    .B(net618),
    .Y(_01961_));
 sky130_fd_sc_hd__xnor2_1 _08004_ (.A(_01960_),
    .B(_01961_),
    .Y(_01962_));
 sky130_fd_sc_hd__nand4_1 _08005_ (.A(net182),
    .B(net427),
    .C(net579),
    .D(net573),
    .Y(_01963_));
 sky130_fd_sc_hd__a22o_1 _08006_ (.A1(net427),
    .A2(net580),
    .B1(net573),
    .B2(net182),
    .X(_01964_));
 sky130_fd_sc_hd__and2_1 _08007_ (.A(net421),
    .B(net588),
    .X(_01965_));
 sky130_fd_sc_hd__a21o_1 _08008_ (.A1(_01963_),
    .A2(_01964_),
    .B1(_01965_),
    .X(_01967_));
 sky130_fd_sc_hd__nand3_1 _08009_ (.A(_01963_),
    .B(_01964_),
    .C(_01965_),
    .Y(_01968_));
 sky130_fd_sc_hd__o21bai_1 _08010_ (.A1(_01792_),
    .A2(_01794_),
    .B1_N(_01793_),
    .Y(_01969_));
 sky130_fd_sc_hd__nand3_2 _08011_ (.A(_01967_),
    .B(_01968_),
    .C(_01969_),
    .Y(_01970_));
 sky130_fd_sc_hd__a21o_1 _08012_ (.A1(_01967_),
    .A2(_01968_),
    .B1(_01969_),
    .X(_01971_));
 sky130_fd_sc_hd__nand3_2 _08013_ (.A(_01962_),
    .B(_01970_),
    .C(_01971_),
    .Y(_01972_));
 sky130_fd_sc_hd__a21o_1 _08014_ (.A1(_01970_),
    .A2(_01971_),
    .B1(_01962_),
    .X(_01973_));
 sky130_fd_sc_hd__and3_1 _08015_ (.A(_01957_),
    .B(_01972_),
    .C(_01973_),
    .X(_01974_));
 sky130_fd_sc_hd__nand3_1 _08016_ (.A(_01957_),
    .B(_01972_),
    .C(_01973_),
    .Y(_01975_));
 sky130_fd_sc_hd__a21oi_1 _08017_ (.A1(_01972_),
    .A2(_01973_),
    .B1(_01957_),
    .Y(_01976_));
 sky130_fd_sc_hd__a211o_1 _08018_ (.A1(_01798_),
    .A2(_01800_),
    .B1(_01974_),
    .C1(_01976_),
    .X(_01978_));
 sky130_fd_sc_hd__o211ai_1 _08019_ (.A1(_01974_),
    .A2(_01976_),
    .B1(_01798_),
    .C1(_01800_),
    .Y(_01979_));
 sky130_fd_sc_hd__and2_1 _08020_ (.A(_01978_),
    .B(_01979_),
    .X(_01980_));
 sky130_fd_sc_hd__nand2_1 _08021_ (.A(_01811_),
    .B(_01814_),
    .Y(_01981_));
 sky130_fd_sc_hd__o21bai_1 _08022_ (.A1(_01819_),
    .A2(_01821_),
    .B1_N(_01820_),
    .Y(_01982_));
 sky130_fd_sc_hd__nand4_1 _08023_ (.A(net209),
    .B(net201),
    .C(net559),
    .D(net552),
    .Y(_01983_));
 sky130_fd_sc_hd__a22o_1 _08024_ (.A1(net201),
    .A2(net559),
    .B1(net552),
    .B2(net209),
    .X(_01984_));
 sky130_fd_sc_hd__a22o_1 _08025_ (.A1(net192),
    .A2(net566),
    .B1(_01983_),
    .B2(_01984_),
    .X(_01985_));
 sky130_fd_sc_hd__nand4_1 _08026_ (.A(net192),
    .B(net566),
    .C(_01983_),
    .D(_01984_),
    .Y(_01986_));
 sky130_fd_sc_hd__and3_1 _08027_ (.A(_01982_),
    .B(_01985_),
    .C(_01986_),
    .X(_01987_));
 sky130_fd_sc_hd__a21o_1 _08028_ (.A1(_01985_),
    .A2(_01986_),
    .B1(_01982_),
    .X(_01989_));
 sky130_fd_sc_hd__and2b_1 _08029_ (.A_N(_01987_),
    .B(_01989_),
    .X(_01990_));
 sky130_fd_sc_hd__xnor2_1 _08030_ (.A(_01981_),
    .B(_01990_),
    .Y(_01991_));
 sky130_fd_sc_hd__nand2_1 _08031_ (.A(net218),
    .B(net538),
    .Y(_01992_));
 sky130_fd_sc_hd__and4_1 _08032_ (.A(net237),
    .B(net229),
    .C(net532),
    .D(net523),
    .X(_01993_));
 sky130_fd_sc_hd__a22oi_1 _08033_ (.A1(net229),
    .A2(net532),
    .B1(net523),
    .B2(net237),
    .Y(_01994_));
 sky130_fd_sc_hd__nor2_1 _08034_ (.A(_01993_),
    .B(_01994_),
    .Y(_01995_));
 sky130_fd_sc_hd__xnor2_1 _08035_ (.A(_01992_),
    .B(_01995_),
    .Y(_01996_));
 sky130_fd_sc_hd__a22oi_1 _08036_ (.A1(net257),
    .A2(net509),
    .B1(net502),
    .B2(net343),
    .Y(_01997_));
 sky130_fd_sc_hd__and4_1 _08037_ (.A(net343),
    .B(net257),
    .C(net509),
    .D(net502),
    .X(_01998_));
 sky130_fd_sc_hd__nor2_1 _08038_ (.A(_01997_),
    .B(_01998_),
    .Y(_02000_));
 sky130_fd_sc_hd__a21boi_1 _08039_ (.A1(_01825_),
    .A2(_01826_),
    .B1_N(_01827_),
    .Y(_02001_));
 sky130_fd_sc_hd__or3_1 _08040_ (.A(_01997_),
    .B(_01998_),
    .C(_02001_),
    .X(_02002_));
 sky130_fd_sc_hd__xnor2_1 _08041_ (.A(_02000_),
    .B(_02001_),
    .Y(_02003_));
 sky130_fd_sc_hd__xnor2_1 _08042_ (.A(_01996_),
    .B(_02003_),
    .Y(_02004_));
 sky130_fd_sc_hd__a21bo_1 _08043_ (.A1(_01823_),
    .A2(_01832_),
    .B1_N(_01831_),
    .X(_02005_));
 sky130_fd_sc_hd__nand2b_1 _08044_ (.A_N(_02004_),
    .B(_02005_),
    .Y(_02006_));
 sky130_fd_sc_hd__xor2_1 _08045_ (.A(_02004_),
    .B(_02005_),
    .X(_02007_));
 sky130_fd_sc_hd__xnor2_1 _08046_ (.A(_01991_),
    .B(_02007_),
    .Y(_02008_));
 sky130_fd_sc_hd__a21bo_1 _08047_ (.A1(_01818_),
    .A2(_01838_),
    .B1_N(_01837_),
    .X(_02009_));
 sky130_fd_sc_hd__and2b_1 _08048_ (.A_N(_02008_),
    .B(_02009_),
    .X(_02011_));
 sky130_fd_sc_hd__xnor2_1 _08049_ (.A(_02008_),
    .B(_02009_),
    .Y(_02012_));
 sky130_fd_sc_hd__xnor2_1 _08050_ (.A(_01980_),
    .B(_02012_),
    .Y(_02013_));
 sky130_fd_sc_hd__a21bo_1 _08051_ (.A1(_01807_),
    .A2(_01842_),
    .B1_N(_01841_),
    .X(_02014_));
 sky130_fd_sc_hd__and2b_1 _08052_ (.A_N(_02013_),
    .B(_02014_),
    .X(_02015_));
 sky130_fd_sc_hd__xnor2_1 _08053_ (.A(_02013_),
    .B(_02014_),
    .Y(_02016_));
 sky130_fd_sc_hd__xor2_1 _08054_ (.A(_01956_),
    .B(_02016_),
    .X(_02017_));
 sky130_fd_sc_hd__a21boi_1 _08055_ (.A1(_01783_),
    .A2(_01847_),
    .B1_N(_01845_),
    .Y(_02018_));
 sky130_fd_sc_hd__and2b_1 _08056_ (.A_N(_02018_),
    .B(_02017_),
    .X(_02019_));
 sky130_fd_sc_hd__xnor2_1 _08057_ (.A(_02017_),
    .B(_02018_),
    .Y(_02020_));
 sky130_fd_sc_hd__xnor2_1 _08058_ (.A(_01917_),
    .B(_02020_),
    .Y(_02022_));
 sky130_fd_sc_hd__a21boi_2 _08059_ (.A1(_01744_),
    .A2(_01851_),
    .B1_N(_01850_),
    .Y(_02023_));
 sky130_fd_sc_hd__or2_1 _08060_ (.A(_02022_),
    .B(_02023_),
    .X(_02024_));
 sky130_fd_sc_hd__xnor2_2 _08061_ (.A(_02022_),
    .B(_02023_),
    .Y(_02025_));
 sky130_fd_sc_hd__xnor2_2 _08062_ (.A(_01870_),
    .B(_02025_),
    .Y(_02026_));
 sky130_fd_sc_hd__a21boi_2 _08063_ (.A1(_01698_),
    .A2(_01855_),
    .B1_N(_01854_),
    .Y(_02027_));
 sky130_fd_sc_hd__or2_1 _08064_ (.A(_02026_),
    .B(_02027_),
    .X(_02028_));
 sky130_fd_sc_hd__xor2_2 _08065_ (.A(_02026_),
    .B(_02027_),
    .X(_02029_));
 sky130_fd_sc_hd__nand2_1 _08066_ (.A(_01868_),
    .B(_02029_),
    .Y(_02030_));
 sky130_fd_sc_hd__xor2_2 _08067_ (.A(_01868_),
    .B(_02029_),
    .X(_02031_));
 sky130_fd_sc_hd__a21boi_2 _08068_ (.A1(_01542_),
    .A2(_01860_),
    .B1_N(_01859_),
    .Y(_02033_));
 sky130_fd_sc_hd__nand2b_1 _08069_ (.A_N(_02033_),
    .B(_02031_),
    .Y(_02034_));
 sky130_fd_sc_hd__xnor2_2 _08070_ (.A(_02031_),
    .B(_02033_),
    .Y(_02035_));
 sky130_fd_sc_hd__or4bb_1 _08071_ (.A(_01692_),
    .B(_01696_),
    .C_N(_01863_),
    .D_N(_01864_),
    .X(_02036_));
 sky130_fd_sc_hd__or3_1 _08072_ (.A(_01059_),
    .B(_01210_),
    .C(_01212_),
    .X(_02037_));
 sky130_fd_sc_hd__o21ba_1 _08073_ (.A1(_01060_),
    .A2(_02037_),
    .B1_N(_01216_),
    .X(_02038_));
 sky130_fd_sc_hd__or3_1 _08074_ (.A(_01692_),
    .B(_01695_),
    .C(_01865_),
    .X(_02039_));
 sky130_fd_sc_hd__a21boi_1 _08075_ (.A1(_01691_),
    .A2(_01863_),
    .B1_N(_01864_),
    .Y(_02040_));
 sky130_fd_sc_hd__o211a_1 _08076_ (.A1(_02036_),
    .A2(_02038_),
    .B1(_02039_),
    .C1(_02040_),
    .X(_02041_));
 sky130_fd_sc_hd__or3_1 _08077_ (.A(_01062_),
    .B(_02036_),
    .C(_02037_),
    .X(_02042_));
 sky130_fd_sc_hd__nand2b_2 _08078_ (.A_N(_02042_),
    .B(_00771_),
    .Y(_02044_));
 sky130_fd_sc_hd__or3b_2 _08079_ (.A(_02042_),
    .B(_05070_),
    .C_N(_00772_),
    .X(_02045_));
 sky130_fd_sc_hd__and3_2 _08080_ (.A(_02041_),
    .B(_02044_),
    .C(_02045_),
    .X(_02046_));
 sky130_fd_sc_hd__inv_2 _08081_ (.A(_02046_),
    .Y(_02047_));
 sky130_fd_sc_hd__xnor2_1 _08082_ (.A(_02035_),
    .B(_02046_),
    .Y(net90));
 sky130_fd_sc_hd__a31o_1 _08083_ (.A1(net602),
    .A2(net248),
    .A3(_01887_),
    .B1(_01886_),
    .X(_02048_));
 sky130_fd_sc_hd__nand2_1 _08084_ (.A(_01914_),
    .B(_01916_),
    .Y(_02049_));
 sky130_fd_sc_hd__a21boi_1 _08085_ (.A1(_01890_),
    .A2(_01910_),
    .B1_N(_01909_),
    .Y(_02050_));
 sky130_fd_sc_hd__o21ai_1 _08086_ (.A1(_01918_),
    .A2(_01954_),
    .B1(_01952_),
    .Y(_02051_));
 sky130_fd_sc_hd__and4_1 _08087_ (.A(net481),
    .B(net473),
    .C(net280),
    .D(net272),
    .X(_02052_));
 sky130_fd_sc_hd__a22oi_1 _08088_ (.A1(net473),
    .A2(net281),
    .B1(net272),
    .B2(net481),
    .Y(_02054_));
 sky130_fd_sc_hd__nor2_1 _08089_ (.A(_02052_),
    .B(_02054_),
    .Y(_02055_));
 sky130_fd_sc_hd__nand2_1 _08090_ (.A(net488),
    .B(net263),
    .Y(_02056_));
 sky130_fd_sc_hd__xnor2_1 _08091_ (.A(_02055_),
    .B(_02056_),
    .Y(_02057_));
 sky130_fd_sc_hd__o21ba_1 _08092_ (.A1(_01874_),
    .A2(_01876_),
    .B1_N(_01873_),
    .X(_02058_));
 sky130_fd_sc_hd__nand2b_1 _08093_ (.A_N(_02058_),
    .B(_02057_),
    .Y(_02059_));
 sky130_fd_sc_hd__xnor2_1 _08094_ (.A(_02057_),
    .B(_02058_),
    .Y(_02060_));
 sky130_fd_sc_hd__nand2_1 _08095_ (.A(net496),
    .B(net252),
    .Y(_02061_));
 sky130_fd_sc_hd__nand3_1 _08096_ (.A(net496),
    .B(net252),
    .C(_02060_),
    .Y(_02062_));
 sky130_fd_sc_hd__xor2_1 _08097_ (.A(_02060_),
    .B(_02061_),
    .X(_02063_));
 sky130_fd_sc_hd__and3_1 _08098_ (.A(_01880_),
    .B(_01883_),
    .C(_02063_),
    .X(_02065_));
 sky130_fd_sc_hd__a21oi_1 _08099_ (.A1(_01880_),
    .A2(_01883_),
    .B1(_02063_),
    .Y(_02066_));
 sky130_fd_sc_hd__nor2_1 _08100_ (.A(_02065_),
    .B(_02066_),
    .Y(_02067_));
 sky130_fd_sc_hd__nand2_1 _08101_ (.A(net517),
    .B(net247),
    .Y(_02068_));
 sky130_fd_sc_hd__xnor2_1 _08102_ (.A(_02067_),
    .B(_02068_),
    .Y(_02069_));
 sky130_fd_sc_hd__a21o_1 _08103_ (.A1(_01924_),
    .A2(_01932_),
    .B1(_01931_),
    .X(_02070_));
 sky130_fd_sc_hd__nand2_1 _08104_ (.A(_01894_),
    .B(_01897_),
    .Y(_02071_));
 sky130_fd_sc_hd__a31o_1 _08105_ (.A1(net442),
    .A2(net317),
    .A3(_01920_),
    .B1(_01919_),
    .X(_02072_));
 sky130_fd_sc_hd__nand4_2 _08106_ (.A(net449),
    .B(net443),
    .C(net309),
    .D(net295),
    .Y(_02073_));
 sky130_fd_sc_hd__a22o_1 _08107_ (.A1(net443),
    .A2(net309),
    .B1(net295),
    .B2(net450),
    .X(_02074_));
 sky130_fd_sc_hd__a22o_1 _08108_ (.A1(net458),
    .A2(net288),
    .B1(_02073_),
    .B2(_02074_),
    .X(_02076_));
 sky130_fd_sc_hd__nand4_2 _08109_ (.A(net458),
    .B(net288),
    .C(_02073_),
    .D(_02074_),
    .Y(_02077_));
 sky130_fd_sc_hd__nand3_2 _08110_ (.A(_02072_),
    .B(_02076_),
    .C(_02077_),
    .Y(_02078_));
 sky130_fd_sc_hd__a21o_1 _08111_ (.A1(_02076_),
    .A2(_02077_),
    .B1(_02072_),
    .X(_02079_));
 sky130_fd_sc_hd__nand3_1 _08112_ (.A(_02071_),
    .B(_02078_),
    .C(_02079_),
    .Y(_02080_));
 sky130_fd_sc_hd__a21o_1 _08113_ (.A1(_02078_),
    .A2(_02079_),
    .B1(_02071_),
    .X(_02081_));
 sky130_fd_sc_hd__and3_1 _08114_ (.A(_02070_),
    .B(_02080_),
    .C(_02081_),
    .X(_02082_));
 sky130_fd_sc_hd__a21oi_1 _08115_ (.A1(_02080_),
    .A2(_02081_),
    .B1(_02070_),
    .Y(_02083_));
 sky130_fd_sc_hd__a211oi_1 _08116_ (.A1(_01898_),
    .A2(_01901_),
    .B1(_02082_),
    .C1(_02083_),
    .Y(_02084_));
 sky130_fd_sc_hd__o211a_1 _08117_ (.A1(_02082_),
    .A2(_02083_),
    .B1(_01898_),
    .C1(_01901_),
    .X(_02085_));
 sky130_fd_sc_hd__nor2_1 _08118_ (.A(_02084_),
    .B(_02085_),
    .Y(_02087_));
 sky130_fd_sc_hd__nor2_1 _08119_ (.A(_01903_),
    .B(_01905_),
    .Y(_02088_));
 sky130_fd_sc_hd__nand2b_1 _08120_ (.A_N(_02088_),
    .B(_02087_),
    .Y(_02089_));
 sky130_fd_sc_hd__xnor2_1 _08121_ (.A(_02087_),
    .B(_02088_),
    .Y(_02090_));
 sky130_fd_sc_hd__xnor2_1 _08122_ (.A(_02069_),
    .B(_02090_),
    .Y(_02091_));
 sky130_fd_sc_hd__nand2b_1 _08123_ (.A_N(_02091_),
    .B(_02051_),
    .Y(_02092_));
 sky130_fd_sc_hd__xor2_1 _08124_ (.A(_02051_),
    .B(_02091_),
    .X(_02093_));
 sky130_fd_sc_hd__xor2_1 _08125_ (.A(_02050_),
    .B(_02093_),
    .X(_02094_));
 sky130_fd_sc_hd__nor2_1 _08126_ (.A(_01948_),
    .B(_01950_),
    .Y(_02095_));
 sky130_fd_sc_hd__and4_1 _08127_ (.A(net463),
    .B(net382),
    .C(net330),
    .D(net323),
    .X(_02096_));
 sky130_fd_sc_hd__a22o_1 _08128_ (.A1(net382),
    .A2(net330),
    .B1(net323),
    .B2(net463),
    .X(_02098_));
 sky130_fd_sc_hd__and2b_1 _08129_ (.A_N(_02096_),
    .B(_02098_),
    .X(_02099_));
 sky130_fd_sc_hd__nand2_1 _08130_ (.A(net543),
    .B(net316),
    .Y(_02100_));
 sky130_fd_sc_hd__xnor2_1 _08131_ (.A(_02099_),
    .B(_02100_),
    .Y(_02101_));
 sky130_fd_sc_hd__nand2_1 _08132_ (.A(net299),
    .B(net339),
    .Y(_02102_));
 sky130_fd_sc_hd__and4_1 _08133_ (.A(net221),
    .B(net177),
    .C(net362),
    .D(net354),
    .X(_02103_));
 sky130_fd_sc_hd__a22oi_2 _08134_ (.A1(net178),
    .A2(net362),
    .B1(net354),
    .B2(net222),
    .Y(_02104_));
 sky130_fd_sc_hd__or3_1 _08135_ (.A(_02102_),
    .B(_02103_),
    .C(_02104_),
    .X(_02105_));
 sky130_fd_sc_hd__o21ai_1 _08136_ (.A1(_02103_),
    .A2(_02104_),
    .B1(_02102_),
    .Y(_02106_));
 sky130_fd_sc_hd__a21bo_1 _08137_ (.A1(_01926_),
    .A2(_01927_),
    .B1_N(_01925_),
    .X(_02107_));
 sky130_fd_sc_hd__and3_1 _08138_ (.A(_02105_),
    .B(_02106_),
    .C(_02107_),
    .X(_02109_));
 sky130_fd_sc_hd__a21o_1 _08139_ (.A1(_02105_),
    .A2(_02106_),
    .B1(_02107_),
    .X(_02110_));
 sky130_fd_sc_hd__and2b_1 _08140_ (.A_N(_02109_),
    .B(_02110_),
    .X(_02111_));
 sky130_fd_sc_hd__xnor2_1 _08141_ (.A(_02101_),
    .B(_02111_),
    .Y(_02112_));
 sky130_fd_sc_hd__nand2_1 _08142_ (.A(_01938_),
    .B(_01941_),
    .Y(_02113_));
 sky130_fd_sc_hd__a31o_1 _08143_ (.A1(net400),
    .A2(net618),
    .A3(_01959_),
    .B1(_01958_),
    .X(_02114_));
 sky130_fd_sc_hd__nand4_1 _08144_ (.A(net392),
    .B(net376),
    .C(net162),
    .D(net618),
    .Y(_02115_));
 sky130_fd_sc_hd__a22o_1 _08145_ (.A1(net376),
    .A2(net162),
    .B1(net619),
    .B2(net392),
    .X(_02116_));
 sky130_fd_sc_hd__a22o_1 _08146_ (.A1(net170),
    .A2(net368),
    .B1(_02115_),
    .B2(_02116_),
    .X(_02117_));
 sky130_fd_sc_hd__nand4_1 _08147_ (.A(net170),
    .B(net369),
    .C(_02115_),
    .D(_02116_),
    .Y(_02118_));
 sky130_fd_sc_hd__nand3_1 _08148_ (.A(_02114_),
    .B(_02117_),
    .C(_02118_),
    .Y(_02120_));
 sky130_fd_sc_hd__a21o_1 _08149_ (.A1(_02117_),
    .A2(_02118_),
    .B1(_02114_),
    .X(_02121_));
 sky130_fd_sc_hd__nand3_1 _08150_ (.A(_02113_),
    .B(_02120_),
    .C(_02121_),
    .Y(_02122_));
 sky130_fd_sc_hd__a21o_1 _08151_ (.A1(_02120_),
    .A2(_02121_),
    .B1(_02113_),
    .X(_02123_));
 sky130_fd_sc_hd__a21bo_1 _08152_ (.A1(_01936_),
    .A2(_01943_),
    .B1_N(_01942_),
    .X(_02124_));
 sky130_fd_sc_hd__and3_1 _08153_ (.A(_02122_),
    .B(_02123_),
    .C(_02124_),
    .X(_02125_));
 sky130_fd_sc_hd__a21oi_1 _08154_ (.A1(_02122_),
    .A2(_02123_),
    .B1(_02124_),
    .Y(_02126_));
 sky130_fd_sc_hd__nor3_1 _08155_ (.A(_02112_),
    .B(_02125_),
    .C(_02126_),
    .Y(_02127_));
 sky130_fd_sc_hd__o21a_1 _08156_ (.A1(_02125_),
    .A2(_02126_),
    .B1(_02112_),
    .X(_02128_));
 sky130_fd_sc_hd__a211o_1 _08157_ (.A1(_01975_),
    .A2(_01978_),
    .B1(_02127_),
    .C1(_02128_),
    .X(_02129_));
 sky130_fd_sc_hd__o211ai_1 _08158_ (.A1(_02127_),
    .A2(_02128_),
    .B1(_01975_),
    .C1(_01978_),
    .Y(_02131_));
 sky130_fd_sc_hd__nand2_1 _08159_ (.A(_02129_),
    .B(_02131_),
    .Y(_02132_));
 sky130_fd_sc_hd__xor2_1 _08160_ (.A(_02095_),
    .B(_02132_),
    .X(_02133_));
 sky130_fd_sc_hd__a21o_1 _08161_ (.A1(_01981_),
    .A2(_01989_),
    .B1(_01987_),
    .X(_02134_));
 sky130_fd_sc_hd__nand2_1 _08162_ (.A(net400),
    .B(net610),
    .Y(_02135_));
 sky130_fd_sc_hd__and4_1 _08163_ (.A(net415),
    .B(net407),
    .C(net594),
    .D(net587),
    .X(_02136_));
 sky130_fd_sc_hd__a22o_1 _08164_ (.A1(net407),
    .A2(net594),
    .B1(net587),
    .B2(net415),
    .X(_02137_));
 sky130_fd_sc_hd__and2b_1 _08165_ (.A_N(_02136_),
    .B(_02137_),
    .X(_02138_));
 sky130_fd_sc_hd__xnor2_1 _08166_ (.A(_02135_),
    .B(_02138_),
    .Y(_02139_));
 sky130_fd_sc_hd__nand2_1 _08167_ (.A(net421),
    .B(net580),
    .Y(_02140_));
 sky130_fd_sc_hd__and4_1 _08168_ (.A(net182),
    .B(net427),
    .C(net573),
    .D(net566),
    .X(_02141_));
 sky130_fd_sc_hd__a22oi_2 _08169_ (.A1(net427),
    .A2(net573),
    .B1(net566),
    .B2(net182),
    .Y(_02142_));
 sky130_fd_sc_hd__or3_1 _08170_ (.A(_02140_),
    .B(_02141_),
    .C(_02142_),
    .X(_02143_));
 sky130_fd_sc_hd__o21ai_1 _08171_ (.A1(_02141_),
    .A2(_02142_),
    .B1(_02140_),
    .Y(_02144_));
 sky130_fd_sc_hd__a21bo_1 _08172_ (.A1(_01964_),
    .A2(_01965_),
    .B1_N(_01963_),
    .X(_02145_));
 sky130_fd_sc_hd__nand3_1 _08173_ (.A(_02143_),
    .B(_02144_),
    .C(_02145_),
    .Y(_02146_));
 sky130_fd_sc_hd__a21o_1 _08174_ (.A1(_02143_),
    .A2(_02144_),
    .B1(_02145_),
    .X(_02147_));
 sky130_fd_sc_hd__nand3_1 _08175_ (.A(_02139_),
    .B(_02146_),
    .C(_02147_),
    .Y(_02148_));
 sky130_fd_sc_hd__a21o_1 _08176_ (.A1(_02146_),
    .A2(_02147_),
    .B1(_02139_),
    .X(_02149_));
 sky130_fd_sc_hd__and3_1 _08177_ (.A(_02134_),
    .B(_02148_),
    .C(_02149_),
    .X(_02150_));
 sky130_fd_sc_hd__a21oi_1 _08178_ (.A1(_02148_),
    .A2(_02149_),
    .B1(_02134_),
    .Y(_02152_));
 sky130_fd_sc_hd__a211oi_2 _08179_ (.A1(_01970_),
    .A2(_01972_),
    .B1(_02150_),
    .C1(_02152_),
    .Y(_02153_));
 sky130_fd_sc_hd__o211a_1 _08180_ (.A1(_02150_),
    .A2(_02152_),
    .B1(_01970_),
    .C1(_01972_),
    .X(_02154_));
 sky130_fd_sc_hd__nor2_1 _08181_ (.A(_02153_),
    .B(_02154_),
    .Y(_02155_));
 sky130_fd_sc_hd__nand2_1 _08182_ (.A(_01983_),
    .B(_01986_),
    .Y(_02156_));
 sky130_fd_sc_hd__o21bai_1 _08183_ (.A1(_01992_),
    .A2(_01994_),
    .B1_N(_01993_),
    .Y(_02157_));
 sky130_fd_sc_hd__nand2_1 _08184_ (.A(net192),
    .B(net559),
    .Y(_02158_));
 sky130_fd_sc_hd__nand4_1 _08185_ (.A(net209),
    .B(net200),
    .C(net552),
    .D(net538),
    .Y(_02159_));
 sky130_fd_sc_hd__a22o_1 _08186_ (.A1(net200),
    .A2(net552),
    .B1(net538),
    .B2(net209),
    .X(_02160_));
 sky130_fd_sc_hd__nand3b_1 _08187_ (.A_N(_02158_),
    .B(_02159_),
    .C(_02160_),
    .Y(_02161_));
 sky130_fd_sc_hd__a21bo_1 _08188_ (.A1(_02159_),
    .A2(_02160_),
    .B1_N(_02158_),
    .X(_02163_));
 sky130_fd_sc_hd__and3_1 _08189_ (.A(_02157_),
    .B(_02161_),
    .C(_02163_),
    .X(_02164_));
 sky130_fd_sc_hd__a21o_1 _08190_ (.A1(_02161_),
    .A2(_02163_),
    .B1(_02157_),
    .X(_02165_));
 sky130_fd_sc_hd__and2b_1 _08191_ (.A_N(_02164_),
    .B(_02165_),
    .X(_02166_));
 sky130_fd_sc_hd__xnor2_1 _08192_ (.A(_02156_),
    .B(_02166_),
    .Y(_02167_));
 sky130_fd_sc_hd__and3_1 _08193_ (.A(net257),
    .B(net502),
    .C(_01650_),
    .X(_02168_));
 sky130_fd_sc_hd__nand2_1 _08194_ (.A(net216),
    .B(net532),
    .Y(_02169_));
 sky130_fd_sc_hd__and4_1 _08195_ (.A(net239),
    .B(net231),
    .C(net523),
    .D(net509),
    .X(_02170_));
 sky130_fd_sc_hd__a22oi_2 _08196_ (.A1(net231),
    .A2(net524),
    .B1(net509),
    .B2(net239),
    .Y(_02171_));
 sky130_fd_sc_hd__or3_1 _08197_ (.A(_02169_),
    .B(_02170_),
    .C(_02171_),
    .X(_02172_));
 sky130_fd_sc_hd__o21ai_1 _08198_ (.A1(_02170_),
    .A2(_02171_),
    .B1(_02169_),
    .Y(_02174_));
 sky130_fd_sc_hd__and3_1 _08199_ (.A(_02168_),
    .B(_02172_),
    .C(_02174_),
    .X(_02175_));
 sky130_fd_sc_hd__a21oi_1 _08200_ (.A1(_02172_),
    .A2(_02174_),
    .B1(_02168_),
    .Y(_02176_));
 sky130_fd_sc_hd__or2_1 _08201_ (.A(_02175_),
    .B(_02176_),
    .X(_02177_));
 sky130_fd_sc_hd__a21bo_1 _08202_ (.A1(_01996_),
    .A2(_02003_),
    .B1_N(_02002_),
    .X(_02178_));
 sky130_fd_sc_hd__and2b_1 _08203_ (.A_N(_02177_),
    .B(_02178_),
    .X(_02179_));
 sky130_fd_sc_hd__xor2_1 _08204_ (.A(_02177_),
    .B(_02178_),
    .X(_02180_));
 sky130_fd_sc_hd__xor2_1 _08205_ (.A(_02167_),
    .B(_02180_),
    .X(_02181_));
 sky130_fd_sc_hd__o21a_1 _08206_ (.A1(_01991_),
    .A2(_02007_),
    .B1(_02006_),
    .X(_02182_));
 sky130_fd_sc_hd__and2b_1 _08207_ (.A_N(_02182_),
    .B(_02181_),
    .X(_02183_));
 sky130_fd_sc_hd__xnor2_1 _08208_ (.A(_02181_),
    .B(_02182_),
    .Y(_02185_));
 sky130_fd_sc_hd__xnor2_1 _08209_ (.A(_02155_),
    .B(_02185_),
    .Y(_02186_));
 sky130_fd_sc_hd__a21oi_1 _08210_ (.A1(_01980_),
    .A2(_02012_),
    .B1(_02011_),
    .Y(_02187_));
 sky130_fd_sc_hd__nor2_1 _08211_ (.A(_02186_),
    .B(_02187_),
    .Y(_02188_));
 sky130_fd_sc_hd__xor2_1 _08212_ (.A(_02186_),
    .B(_02187_),
    .X(_02189_));
 sky130_fd_sc_hd__xor2_1 _08213_ (.A(_02133_),
    .B(_02189_),
    .X(_02190_));
 sky130_fd_sc_hd__a21oi_1 _08214_ (.A1(_01956_),
    .A2(_02016_),
    .B1(_02015_),
    .Y(_02191_));
 sky130_fd_sc_hd__and2b_1 _08215_ (.A_N(_02191_),
    .B(_02190_),
    .X(_02192_));
 sky130_fd_sc_hd__xnor2_1 _08216_ (.A(_02190_),
    .B(_02191_),
    .Y(_02193_));
 sky130_fd_sc_hd__xnor2_1 _08217_ (.A(_02094_),
    .B(_02193_),
    .Y(_02194_));
 sky130_fd_sc_hd__a21oi_1 _08218_ (.A1(_01917_),
    .A2(_02020_),
    .B1(_02019_),
    .Y(_02196_));
 sky130_fd_sc_hd__nor2_1 _08219_ (.A(_02194_),
    .B(_02196_),
    .Y(_02197_));
 sky130_fd_sc_hd__nand2_1 _08220_ (.A(_02194_),
    .B(_02196_),
    .Y(_02198_));
 sky130_fd_sc_hd__xnor2_1 _08221_ (.A(_02194_),
    .B(_02196_),
    .Y(_02199_));
 sky130_fd_sc_hd__xnor2_1 _08222_ (.A(_02049_),
    .B(_02199_),
    .Y(_02200_));
 sky130_fd_sc_hd__o21a_1 _08223_ (.A1(_01870_),
    .A2(_02025_),
    .B1(_02024_),
    .X(_02201_));
 sky130_fd_sc_hd__nand2b_1 _08224_ (.A_N(_02201_),
    .B(_02200_),
    .Y(_02202_));
 sky130_fd_sc_hd__xnor2_1 _08225_ (.A(_02200_),
    .B(_02201_),
    .Y(_02203_));
 sky130_fd_sc_hd__xnor2_1 _08226_ (.A(_02048_),
    .B(_02203_),
    .Y(_02204_));
 sky130_fd_sc_hd__a21o_1 _08227_ (.A1(_02028_),
    .A2(_02030_),
    .B1(_02204_),
    .X(_02205_));
 sky130_fd_sc_hd__inv_2 _08228_ (.A(_02205_),
    .Y(_02207_));
 sky130_fd_sc_hd__and3_1 _08229_ (.A(_02028_),
    .B(_02030_),
    .C(_02204_),
    .X(_02208_));
 sky130_fd_sc_hd__nor2_1 _08230_ (.A(_02207_),
    .B(_02208_),
    .Y(_02209_));
 sky130_fd_sc_hd__a21bo_1 _08231_ (.A1(_02035_),
    .A2(_02047_),
    .B1_N(_02034_),
    .X(_02210_));
 sky130_fd_sc_hd__xor2_1 _08232_ (.A(_02209_),
    .B(_02210_),
    .X(net91));
 sky130_fd_sc_hd__a31o_1 _08233_ (.A1(net517),
    .A2(net247),
    .A3(_02067_),
    .B1(_02066_),
    .X(_02211_));
 sky130_fd_sc_hd__o21ai_1 _08234_ (.A1(_02050_),
    .A2(_02093_),
    .B1(_02092_),
    .Y(_02212_));
 sky130_fd_sc_hd__a21boi_1 _08235_ (.A1(_02069_),
    .A2(_02090_),
    .B1_N(_02089_),
    .Y(_02213_));
 sky130_fd_sc_hd__o21ai_1 _08236_ (.A1(_02095_),
    .A2(_02132_),
    .B1(_02129_),
    .Y(_02214_));
 sky130_fd_sc_hd__and4_1 _08237_ (.A(net473),
    .B(net458),
    .C(net280),
    .D(net272),
    .X(_02215_));
 sky130_fd_sc_hd__a22oi_1 _08238_ (.A1(net458),
    .A2(net280),
    .B1(net272),
    .B2(net473),
    .Y(_02217_));
 sky130_fd_sc_hd__nor2_1 _08239_ (.A(_02215_),
    .B(_02217_),
    .Y(_02218_));
 sky130_fd_sc_hd__nand2_1 _08240_ (.A(net481),
    .B(net263),
    .Y(_02219_));
 sky130_fd_sc_hd__xnor2_1 _08241_ (.A(_02218_),
    .B(_02219_),
    .Y(_02220_));
 sky130_fd_sc_hd__o21ba_1 _08242_ (.A1(_02054_),
    .A2(_02056_),
    .B1_N(_02052_),
    .X(_02221_));
 sky130_fd_sc_hd__nand2b_1 _08243_ (.A_N(_02221_),
    .B(_02220_),
    .Y(_02222_));
 sky130_fd_sc_hd__xnor2_1 _08244_ (.A(_02220_),
    .B(_02221_),
    .Y(_02223_));
 sky130_fd_sc_hd__nand2_1 _08245_ (.A(net488),
    .B(net252),
    .Y(_02224_));
 sky130_fd_sc_hd__nand3_1 _08246_ (.A(net488),
    .B(net252),
    .C(_02223_),
    .Y(_02225_));
 sky130_fd_sc_hd__xor2_1 _08247_ (.A(_02223_),
    .B(_02224_),
    .X(_02226_));
 sky130_fd_sc_hd__and3_1 _08248_ (.A(_02059_),
    .B(_02062_),
    .C(_02226_),
    .X(_02228_));
 sky130_fd_sc_hd__a21oi_1 _08249_ (.A1(_02059_),
    .A2(_02062_),
    .B1(_02226_),
    .Y(_02229_));
 sky130_fd_sc_hd__nor2_1 _08250_ (.A(_02228_),
    .B(_02229_),
    .Y(_02230_));
 sky130_fd_sc_hd__nand2_1 _08251_ (.A(net496),
    .B(net247),
    .Y(_02231_));
 sky130_fd_sc_hd__xnor2_1 _08252_ (.A(_02230_),
    .B(_02231_),
    .Y(_02232_));
 sky130_fd_sc_hd__a21o_1 _08253_ (.A1(_02101_),
    .A2(_02110_),
    .B1(_02109_),
    .X(_02233_));
 sky130_fd_sc_hd__nand2_1 _08254_ (.A(_02073_),
    .B(_02077_),
    .Y(_02234_));
 sky130_fd_sc_hd__a31o_1 _08255_ (.A1(net543),
    .A2(net316),
    .A3(_02098_),
    .B1(_02096_),
    .X(_02235_));
 sky130_fd_sc_hd__nand4_2 _08256_ (.A(net543),
    .B(net442),
    .C(net308),
    .D(net294),
    .Y(_02236_));
 sky130_fd_sc_hd__a22o_1 _08257_ (.A1(net543),
    .A2(net308),
    .B1(net294),
    .B2(net442),
    .X(_02237_));
 sky130_fd_sc_hd__a22o_1 _08258_ (.A1(net449),
    .A2(net287),
    .B1(_02236_),
    .B2(_02237_),
    .X(_02239_));
 sky130_fd_sc_hd__nand4_2 _08259_ (.A(net449),
    .B(net287),
    .C(_02236_),
    .D(_02237_),
    .Y(_02240_));
 sky130_fd_sc_hd__nand3_2 _08260_ (.A(_02235_),
    .B(_02239_),
    .C(_02240_),
    .Y(_02241_));
 sky130_fd_sc_hd__a21o_1 _08261_ (.A1(_02239_),
    .A2(_02240_),
    .B1(_02235_),
    .X(_02242_));
 sky130_fd_sc_hd__nand3_2 _08262_ (.A(_02234_),
    .B(_02241_),
    .C(_02242_),
    .Y(_02243_));
 sky130_fd_sc_hd__a21o_1 _08263_ (.A1(_02241_),
    .A2(_02242_),
    .B1(_02234_),
    .X(_02244_));
 sky130_fd_sc_hd__and3_1 _08264_ (.A(_02233_),
    .B(_02243_),
    .C(_02244_),
    .X(_02245_));
 sky130_fd_sc_hd__a21oi_1 _08265_ (.A1(_02243_),
    .A2(_02244_),
    .B1(_02233_),
    .Y(_02246_));
 sky130_fd_sc_hd__a211oi_1 _08266_ (.A1(_02078_),
    .A2(_02080_),
    .B1(_02245_),
    .C1(_02246_),
    .Y(_02247_));
 sky130_fd_sc_hd__o211a_1 _08267_ (.A1(_02245_),
    .A2(_02246_),
    .B1(_02078_),
    .C1(_02080_),
    .X(_02248_));
 sky130_fd_sc_hd__nor2_1 _08268_ (.A(_02247_),
    .B(_02248_),
    .Y(_02250_));
 sky130_fd_sc_hd__nor2_1 _08269_ (.A(_02082_),
    .B(_02084_),
    .Y(_02251_));
 sky130_fd_sc_hd__nand2b_1 _08270_ (.A_N(_02251_),
    .B(_02250_),
    .Y(_02252_));
 sky130_fd_sc_hd__xnor2_1 _08271_ (.A(_02250_),
    .B(_02251_),
    .Y(_02253_));
 sky130_fd_sc_hd__xnor2_1 _08272_ (.A(_02232_),
    .B(_02253_),
    .Y(_02254_));
 sky130_fd_sc_hd__nand2b_1 _08273_ (.A_N(_02254_),
    .B(_02214_),
    .Y(_02255_));
 sky130_fd_sc_hd__xor2_1 _08274_ (.A(_02214_),
    .B(_02254_),
    .X(_02256_));
 sky130_fd_sc_hd__xor2_1 _08275_ (.A(_02213_),
    .B(_02256_),
    .X(_02257_));
 sky130_fd_sc_hd__nor2_1 _08276_ (.A(_02125_),
    .B(_02127_),
    .Y(_02258_));
 sky130_fd_sc_hd__and4_1 _08277_ (.A(net382),
    .B(net298),
    .C(net330),
    .D(net323),
    .X(_02259_));
 sky130_fd_sc_hd__a22o_1 _08278_ (.A1(net298),
    .A2(net330),
    .B1(net323),
    .B2(net382),
    .X(_02261_));
 sky130_fd_sc_hd__and2b_1 _08279_ (.A_N(_02259_),
    .B(_02261_),
    .X(_02262_));
 sky130_fd_sc_hd__nand2_1 _08280_ (.A(net463),
    .B(net316),
    .Y(_02263_));
 sky130_fd_sc_hd__xnor2_1 _08281_ (.A(_02262_),
    .B(_02263_),
    .Y(_02264_));
 sky130_fd_sc_hd__nand2_1 _08282_ (.A(net221),
    .B(net339),
    .Y(_02265_));
 sky130_fd_sc_hd__and4_1 _08283_ (.A(net177),
    .B(net169),
    .C(net362),
    .D(net354),
    .X(_02266_));
 sky130_fd_sc_hd__a22oi_2 _08284_ (.A1(net170),
    .A2(net362),
    .B1(net354),
    .B2(net178),
    .Y(_02267_));
 sky130_fd_sc_hd__or3_1 _08285_ (.A(_02265_),
    .B(_02266_),
    .C(_02267_),
    .X(_02268_));
 sky130_fd_sc_hd__o21ai_1 _08286_ (.A1(_02266_),
    .A2(_02267_),
    .B1(_02265_),
    .Y(_02269_));
 sky130_fd_sc_hd__o21bai_1 _08287_ (.A1(_02102_),
    .A2(_02104_),
    .B1_N(_02103_),
    .Y(_02270_));
 sky130_fd_sc_hd__and3_1 _08288_ (.A(_02268_),
    .B(_02269_),
    .C(_02270_),
    .X(_02272_));
 sky130_fd_sc_hd__a21o_1 _08289_ (.A1(_02268_),
    .A2(_02269_),
    .B1(_02270_),
    .X(_02273_));
 sky130_fd_sc_hd__and2b_1 _08290_ (.A_N(_02272_),
    .B(_02273_),
    .X(_02274_));
 sky130_fd_sc_hd__xnor2_1 _08291_ (.A(_02264_),
    .B(_02274_),
    .Y(_02275_));
 sky130_fd_sc_hd__nand2_1 _08292_ (.A(_02115_),
    .B(_02118_),
    .Y(_02276_));
 sky130_fd_sc_hd__a31o_1 _08293_ (.A1(net400),
    .A2(net611),
    .A3(_02137_),
    .B1(_02136_),
    .X(_02277_));
 sky130_fd_sc_hd__nand4_1 _08294_ (.A(net391),
    .B(net375),
    .C(net618),
    .D(net610),
    .Y(_02278_));
 sky130_fd_sc_hd__a22o_1 _08295_ (.A1(net376),
    .A2(net619),
    .B1(net610),
    .B2(net392),
    .X(_02279_));
 sky130_fd_sc_hd__a22o_1 _08296_ (.A1(net162),
    .A2(net369),
    .B1(_02278_),
    .B2(_02279_),
    .X(_02280_));
 sky130_fd_sc_hd__nand4_1 _08297_ (.A(net162),
    .B(net369),
    .C(_02278_),
    .D(_02279_),
    .Y(_02281_));
 sky130_fd_sc_hd__nand3_1 _08298_ (.A(_02277_),
    .B(_02280_),
    .C(_02281_),
    .Y(_02283_));
 sky130_fd_sc_hd__a21o_1 _08299_ (.A1(_02280_),
    .A2(_02281_),
    .B1(_02277_),
    .X(_02284_));
 sky130_fd_sc_hd__nand3_1 _08300_ (.A(_02276_),
    .B(_02283_),
    .C(_02284_),
    .Y(_02285_));
 sky130_fd_sc_hd__a21o_1 _08301_ (.A1(_02283_),
    .A2(_02284_),
    .B1(_02276_),
    .X(_02286_));
 sky130_fd_sc_hd__a21bo_1 _08302_ (.A1(_02113_),
    .A2(_02121_),
    .B1_N(_02120_),
    .X(_02287_));
 sky130_fd_sc_hd__and3_1 _08303_ (.A(_02285_),
    .B(_02286_),
    .C(_02287_),
    .X(_02288_));
 sky130_fd_sc_hd__a21oi_1 _08304_ (.A1(_02285_),
    .A2(_02286_),
    .B1(_02287_),
    .Y(_02289_));
 sky130_fd_sc_hd__or3_1 _08305_ (.A(_02275_),
    .B(_02288_),
    .C(_02289_),
    .X(_02290_));
 sky130_fd_sc_hd__o21ai_1 _08306_ (.A1(_02288_),
    .A2(_02289_),
    .B1(_02275_),
    .Y(_02291_));
 sky130_fd_sc_hd__o211ai_1 _08307_ (.A1(_02150_),
    .A2(_02153_),
    .B1(_02290_),
    .C1(_02291_),
    .Y(_02292_));
 sky130_fd_sc_hd__a211o_1 _08308_ (.A1(_02290_),
    .A2(_02291_),
    .B1(_02150_),
    .C1(_02153_),
    .X(_02294_));
 sky130_fd_sc_hd__nand2_1 _08309_ (.A(_02292_),
    .B(_02294_),
    .Y(_02295_));
 sky130_fd_sc_hd__xor2_1 _08310_ (.A(_02258_),
    .B(_02295_),
    .X(_02296_));
 sky130_fd_sc_hd__nand2_1 _08311_ (.A(_02146_),
    .B(_02148_),
    .Y(_02297_));
 sky130_fd_sc_hd__a21o_1 _08312_ (.A1(_02156_),
    .A2(_02165_),
    .B1(_02164_),
    .X(_02298_));
 sky130_fd_sc_hd__nand2_1 _08313_ (.A(net399),
    .B(net594),
    .Y(_02299_));
 sky130_fd_sc_hd__and4_1 _08314_ (.A(net414),
    .B(net406),
    .C(net587),
    .D(net579),
    .X(_02300_));
 sky130_fd_sc_hd__a22o_1 _08315_ (.A1(net406),
    .A2(net587),
    .B1(net579),
    .B2(net414),
    .X(_02301_));
 sky130_fd_sc_hd__and2b_1 _08316_ (.A_N(_02300_),
    .B(_02301_),
    .X(_02302_));
 sky130_fd_sc_hd__xnor2_1 _08317_ (.A(_02299_),
    .B(_02302_),
    .Y(_02303_));
 sky130_fd_sc_hd__nand2_1 _08318_ (.A(net421),
    .B(net574),
    .Y(_02305_));
 sky130_fd_sc_hd__and4_1 _08319_ (.A(net182),
    .B(net427),
    .C(net566),
    .D(net559),
    .X(_02306_));
 sky130_fd_sc_hd__a22oi_2 _08320_ (.A1(net427),
    .A2(net566),
    .B1(net559),
    .B2(net182),
    .Y(_02307_));
 sky130_fd_sc_hd__or3_1 _08321_ (.A(_02305_),
    .B(_02306_),
    .C(_02307_),
    .X(_02308_));
 sky130_fd_sc_hd__o21ai_1 _08322_ (.A1(_02306_),
    .A2(_02307_),
    .B1(_02305_),
    .Y(_02309_));
 sky130_fd_sc_hd__o21bai_1 _08323_ (.A1(_02140_),
    .A2(_02142_),
    .B1_N(_02141_),
    .Y(_02310_));
 sky130_fd_sc_hd__nand3_1 _08324_ (.A(_02308_),
    .B(_02309_),
    .C(_02310_),
    .Y(_02311_));
 sky130_fd_sc_hd__a21o_1 _08325_ (.A1(_02308_),
    .A2(_02309_),
    .B1(_02310_),
    .X(_02312_));
 sky130_fd_sc_hd__nand3_1 _08326_ (.A(_02303_),
    .B(_02311_),
    .C(_02312_),
    .Y(_02313_));
 sky130_fd_sc_hd__a21o_1 _08327_ (.A1(_02311_),
    .A2(_02312_),
    .B1(_02303_),
    .X(_02314_));
 sky130_fd_sc_hd__nand3_2 _08328_ (.A(_02298_),
    .B(_02313_),
    .C(_02314_),
    .Y(_02316_));
 sky130_fd_sc_hd__a21o_1 _08329_ (.A1(_02313_),
    .A2(_02314_),
    .B1(_02298_),
    .X(_02317_));
 sky130_fd_sc_hd__nand3_1 _08330_ (.A(_02297_),
    .B(_02316_),
    .C(_02317_),
    .Y(_02318_));
 sky130_fd_sc_hd__a21o_1 _08331_ (.A1(_02316_),
    .A2(_02317_),
    .B1(_02297_),
    .X(_02319_));
 sky130_fd_sc_hd__and2_1 _08332_ (.A(_02318_),
    .B(_02319_),
    .X(_02320_));
 sky130_fd_sc_hd__nand2_1 _08333_ (.A(_02159_),
    .B(_02161_),
    .Y(_02321_));
 sky130_fd_sc_hd__o21bai_1 _08334_ (.A1(_02169_),
    .A2(_02171_),
    .B1_N(_02170_),
    .Y(_02322_));
 sky130_fd_sc_hd__nand2_1 _08335_ (.A(net192),
    .B(net552),
    .Y(_02323_));
 sky130_fd_sc_hd__nand4_1 _08336_ (.A(net211),
    .B(net200),
    .C(net542),
    .D(net532),
    .Y(_02324_));
 sky130_fd_sc_hd__a22o_1 _08337_ (.A1(net200),
    .A2(net542),
    .B1(net533),
    .B2(net211),
    .X(_02325_));
 sky130_fd_sc_hd__nand3b_1 _08338_ (.A_N(_02323_),
    .B(_02324_),
    .C(_02325_),
    .Y(_02327_));
 sky130_fd_sc_hd__a21bo_1 _08339_ (.A1(_02324_),
    .A2(_02325_),
    .B1_N(_02323_),
    .X(_02328_));
 sky130_fd_sc_hd__nand3_1 _08340_ (.A(_02322_),
    .B(_02327_),
    .C(_02328_),
    .Y(_02329_));
 sky130_fd_sc_hd__a21o_1 _08341_ (.A1(_02327_),
    .A2(_02328_),
    .B1(_02322_),
    .X(_02330_));
 sky130_fd_sc_hd__nand3_1 _08342_ (.A(_02321_),
    .B(_02329_),
    .C(_02330_),
    .Y(_02331_));
 sky130_fd_sc_hd__a21o_1 _08343_ (.A1(_02329_),
    .A2(_02330_),
    .B1(_02321_),
    .X(_02332_));
 sky130_fd_sc_hd__and2_1 _08344_ (.A(_02331_),
    .B(_02332_),
    .X(_02333_));
 sky130_fd_sc_hd__nand2_1 _08345_ (.A(net216),
    .B(net524),
    .Y(_02334_));
 sky130_fd_sc_hd__and4_1 _08346_ (.A(net239),
    .B(net231),
    .C(net509),
    .D(net502),
    .X(_02335_));
 sky130_fd_sc_hd__a22o_1 _08347_ (.A1(net231),
    .A2(net509),
    .B1(net502),
    .B2(net239),
    .X(_02336_));
 sky130_fd_sc_hd__and2b_1 _08348_ (.A_N(_02335_),
    .B(_02336_),
    .X(_02338_));
 sky130_fd_sc_hd__xnor2_1 _08349_ (.A(_02334_),
    .B(_02338_),
    .Y(_02339_));
 sky130_fd_sc_hd__o21a_1 _08350_ (.A1(_01998_),
    .A2(_02175_),
    .B1(_02339_),
    .X(_02340_));
 sky130_fd_sc_hd__or3_1 _08351_ (.A(_01998_),
    .B(_02175_),
    .C(_02339_),
    .X(_02341_));
 sky130_fd_sc_hd__and2b_1 _08352_ (.A_N(_02340_),
    .B(_02341_),
    .X(_02342_));
 sky130_fd_sc_hd__xnor2_1 _08353_ (.A(_02333_),
    .B(_02342_),
    .Y(_02343_));
 sky130_fd_sc_hd__o21ba_1 _08354_ (.A1(_02167_),
    .A2(_02180_),
    .B1_N(_02179_),
    .X(_02344_));
 sky130_fd_sc_hd__nor2_1 _08355_ (.A(_02343_),
    .B(_02344_),
    .Y(_02345_));
 sky130_fd_sc_hd__xor2_1 _08356_ (.A(_02343_),
    .B(_02344_),
    .X(_02346_));
 sky130_fd_sc_hd__xnor2_1 _08357_ (.A(_02320_),
    .B(_02346_),
    .Y(_02347_));
 sky130_fd_sc_hd__a21oi_1 _08358_ (.A1(_02155_),
    .A2(_02185_),
    .B1(_02183_),
    .Y(_02349_));
 sky130_fd_sc_hd__nor2_1 _08359_ (.A(_02347_),
    .B(_02349_),
    .Y(_02350_));
 sky130_fd_sc_hd__xor2_1 _08360_ (.A(_02347_),
    .B(_02349_),
    .X(_02351_));
 sky130_fd_sc_hd__xor2_1 _08361_ (.A(_02296_),
    .B(_02351_),
    .X(_02352_));
 sky130_fd_sc_hd__a21oi_1 _08362_ (.A1(_02133_),
    .A2(_02189_),
    .B1(_02188_),
    .Y(_02353_));
 sky130_fd_sc_hd__and2b_1 _08363_ (.A_N(_02353_),
    .B(_02352_),
    .X(_02354_));
 sky130_fd_sc_hd__xnor2_1 _08364_ (.A(_02352_),
    .B(_02353_),
    .Y(_02355_));
 sky130_fd_sc_hd__xnor2_1 _08365_ (.A(_02257_),
    .B(_02355_),
    .Y(_02356_));
 sky130_fd_sc_hd__a21oi_1 _08366_ (.A1(_02094_),
    .A2(_02193_),
    .B1(_02192_),
    .Y(_02357_));
 sky130_fd_sc_hd__nor2_1 _08367_ (.A(_02356_),
    .B(_02357_),
    .Y(_02358_));
 sky130_fd_sc_hd__nand2_1 _08368_ (.A(_02356_),
    .B(_02357_),
    .Y(_02360_));
 sky130_fd_sc_hd__xnor2_1 _08369_ (.A(_02356_),
    .B(_02357_),
    .Y(_02361_));
 sky130_fd_sc_hd__xnor2_1 _08370_ (.A(_02212_),
    .B(_02361_),
    .Y(_02362_));
 sky130_fd_sc_hd__a21oi_1 _08371_ (.A1(_02049_),
    .A2(_02198_),
    .B1(_02197_),
    .Y(_02363_));
 sky130_fd_sc_hd__nand2b_1 _08372_ (.A_N(_02363_),
    .B(_02362_),
    .Y(_02364_));
 sky130_fd_sc_hd__xnor2_1 _08373_ (.A(_02362_),
    .B(_02363_),
    .Y(_02365_));
 sky130_fd_sc_hd__nand2_1 _08374_ (.A(_02211_),
    .B(_02365_),
    .Y(_02366_));
 sky130_fd_sc_hd__xnor2_1 _08375_ (.A(_02211_),
    .B(_02365_),
    .Y(_02367_));
 sky130_fd_sc_hd__a21boi_1 _08376_ (.A1(_02048_),
    .A2(_02203_),
    .B1_N(_02202_),
    .Y(_02368_));
 sky130_fd_sc_hd__or2_1 _08377_ (.A(_02367_),
    .B(_02368_),
    .X(_02369_));
 sky130_fd_sc_hd__nand2_1 _08378_ (.A(_02367_),
    .B(_02368_),
    .Y(_02371_));
 sky130_fd_sc_hd__xnor2_1 _08379_ (.A(_02367_),
    .B(_02368_),
    .Y(_02372_));
 sky130_fd_sc_hd__a21o_1 _08380_ (.A1(_02034_),
    .A2(_02205_),
    .B1(_02208_),
    .X(_02373_));
 sky130_fd_sc_hd__nand2_1 _08381_ (.A(_02035_),
    .B(_02209_),
    .Y(_02374_));
 sky130_fd_sc_hd__o21ai_1 _08382_ (.A1(_02046_),
    .A2(_02374_),
    .B1(_02373_),
    .Y(_02375_));
 sky130_fd_sc_hd__xnor2_1 _08383_ (.A(_02372_),
    .B(_02375_),
    .Y(net92));
 sky130_fd_sc_hd__a31o_1 _08384_ (.A1(net496),
    .A2(net247),
    .A3(_02230_),
    .B1(_02229_),
    .X(_02376_));
 sky130_fd_sc_hd__o21ai_1 _08385_ (.A1(_02213_),
    .A2(_02256_),
    .B1(_02255_),
    .Y(_02377_));
 sky130_fd_sc_hd__inv_2 _08386_ (.A(_02377_),
    .Y(_02378_));
 sky130_fd_sc_hd__a21boi_1 _08387_ (.A1(_02232_),
    .A2(_02253_),
    .B1_N(_02252_),
    .Y(_02379_));
 sky130_fd_sc_hd__o21ai_1 _08388_ (.A1(_02258_),
    .A2(_02295_),
    .B1(_02292_),
    .Y(_02381_));
 sky130_fd_sc_hd__and4_1 _08389_ (.A(net458),
    .B(net450),
    .C(net280),
    .D(net273),
    .X(_02382_));
 sky130_fd_sc_hd__a22oi_1 _08390_ (.A1(net450),
    .A2(net280),
    .B1(net273),
    .B2(net458),
    .Y(_02383_));
 sky130_fd_sc_hd__o2bb2a_1 _08391_ (.A1_N(net473),
    .A2_N(net263),
    .B1(_02382_),
    .B2(_02383_),
    .X(_02384_));
 sky130_fd_sc_hd__and4bb_1 _08392_ (.A_N(_02382_),
    .B_N(_02383_),
    .C(net473),
    .D(net263),
    .X(_02385_));
 sky130_fd_sc_hd__nor2_1 _08393_ (.A(_02384_),
    .B(_02385_),
    .Y(_02386_));
 sky130_fd_sc_hd__o21ba_1 _08394_ (.A1(_02217_),
    .A2(_02219_),
    .B1_N(_02215_),
    .X(_02387_));
 sky130_fd_sc_hd__or3_1 _08395_ (.A(_02384_),
    .B(_02385_),
    .C(_02387_),
    .X(_02388_));
 sky130_fd_sc_hd__xnor2_1 _08396_ (.A(_02386_),
    .B(_02387_),
    .Y(_02389_));
 sky130_fd_sc_hd__nand2_1 _08397_ (.A(net481),
    .B(net252),
    .Y(_02390_));
 sky130_fd_sc_hd__nand3_1 _08398_ (.A(net481),
    .B(net252),
    .C(_02389_),
    .Y(_02392_));
 sky130_fd_sc_hd__xor2_1 _08399_ (.A(_02389_),
    .B(_02390_),
    .X(_02393_));
 sky130_fd_sc_hd__and3_1 _08400_ (.A(_02222_),
    .B(_02225_),
    .C(_02393_),
    .X(_02394_));
 sky130_fd_sc_hd__a21oi_1 _08401_ (.A1(_02222_),
    .A2(_02225_),
    .B1(_02393_),
    .Y(_02395_));
 sky130_fd_sc_hd__nor2_1 _08402_ (.A(_02394_),
    .B(_02395_),
    .Y(_02396_));
 sky130_fd_sc_hd__nand2_1 _08403_ (.A(net488),
    .B(net247),
    .Y(_02397_));
 sky130_fd_sc_hd__xnor2_1 _08404_ (.A(_02396_),
    .B(_02397_),
    .Y(_02398_));
 sky130_fd_sc_hd__a21o_1 _08405_ (.A1(_02264_),
    .A2(_02273_),
    .B1(_02272_),
    .X(_02399_));
 sky130_fd_sc_hd__nand2_1 _08406_ (.A(_02236_),
    .B(_02240_),
    .Y(_02400_));
 sky130_fd_sc_hd__a31o_1 _08407_ (.A1(net463),
    .A2(net316),
    .A3(_02261_),
    .B1(_02259_),
    .X(_02401_));
 sky130_fd_sc_hd__nand4_2 _08408_ (.A(net543),
    .B(net463),
    .C(net308),
    .D(net294),
    .Y(_02403_));
 sky130_fd_sc_hd__a22o_1 _08409_ (.A1(net463),
    .A2(net308),
    .B1(net294),
    .B2(net543),
    .X(_02404_));
 sky130_fd_sc_hd__a22o_1 _08410_ (.A1(net442),
    .A2(net287),
    .B1(_02403_),
    .B2(_02404_),
    .X(_02405_));
 sky130_fd_sc_hd__nand4_2 _08411_ (.A(net442),
    .B(net287),
    .C(_02403_),
    .D(_02404_),
    .Y(_02406_));
 sky130_fd_sc_hd__nand3_2 _08412_ (.A(_02401_),
    .B(_02405_),
    .C(_02406_),
    .Y(_02407_));
 sky130_fd_sc_hd__a21o_1 _08413_ (.A1(_02405_),
    .A2(_02406_),
    .B1(_02401_),
    .X(_02408_));
 sky130_fd_sc_hd__nand3_2 _08414_ (.A(_02400_),
    .B(_02407_),
    .C(_02408_),
    .Y(_02409_));
 sky130_fd_sc_hd__a21o_1 _08415_ (.A1(_02407_),
    .A2(_02408_),
    .B1(_02400_),
    .X(_02410_));
 sky130_fd_sc_hd__and3_1 _08416_ (.A(_02399_),
    .B(_02409_),
    .C(_02410_),
    .X(_02411_));
 sky130_fd_sc_hd__a21oi_1 _08417_ (.A1(_02409_),
    .A2(_02410_),
    .B1(_02399_),
    .Y(_02412_));
 sky130_fd_sc_hd__a211oi_1 _08418_ (.A1(_02241_),
    .A2(_02243_),
    .B1(_02411_),
    .C1(_02412_),
    .Y(_02414_));
 sky130_fd_sc_hd__a211o_1 _08419_ (.A1(_02241_),
    .A2(_02243_),
    .B1(_02411_),
    .C1(_02412_),
    .X(_02415_));
 sky130_fd_sc_hd__o211ai_1 _08420_ (.A1(_02411_),
    .A2(_02412_),
    .B1(_02241_),
    .C1(_02243_),
    .Y(_02416_));
 sky130_fd_sc_hd__o211ai_1 _08421_ (.A1(_02245_),
    .A2(_02247_),
    .B1(_02415_),
    .C1(_02416_),
    .Y(_02417_));
 sky130_fd_sc_hd__a211o_1 _08422_ (.A1(_02415_),
    .A2(_02416_),
    .B1(_02245_),
    .C1(_02247_),
    .X(_02418_));
 sky130_fd_sc_hd__nand2_1 _08423_ (.A(_02417_),
    .B(_02418_),
    .Y(_02419_));
 sky130_fd_sc_hd__xor2_1 _08424_ (.A(_02398_),
    .B(_02419_),
    .X(_02420_));
 sky130_fd_sc_hd__nand2b_1 _08425_ (.A_N(_02420_),
    .B(_02381_),
    .Y(_02421_));
 sky130_fd_sc_hd__xor2_1 _08426_ (.A(_02381_),
    .B(_02420_),
    .X(_02422_));
 sky130_fd_sc_hd__xor2_1 _08427_ (.A(_02379_),
    .B(_02422_),
    .X(_02423_));
 sky130_fd_sc_hd__and2b_1 _08428_ (.A_N(_02288_),
    .B(_02290_),
    .X(_02425_));
 sky130_fd_sc_hd__and4_1 _08429_ (.A(net298),
    .B(net221),
    .C(net330),
    .D(net323),
    .X(_02426_));
 sky130_fd_sc_hd__a22o_1 _08430_ (.A1(net221),
    .A2(net330),
    .B1(net323),
    .B2(net298),
    .X(_02427_));
 sky130_fd_sc_hd__and2b_1 _08431_ (.A_N(_02426_),
    .B(_02427_),
    .X(_02428_));
 sky130_fd_sc_hd__nand2_1 _08432_ (.A(net382),
    .B(net316),
    .Y(_02429_));
 sky130_fd_sc_hd__xnor2_1 _08433_ (.A(_02428_),
    .B(_02429_),
    .Y(_02430_));
 sky130_fd_sc_hd__nand2_1 _08434_ (.A(net177),
    .B(net339),
    .Y(_02431_));
 sky130_fd_sc_hd__and4_1 _08435_ (.A(net169),
    .B(net161),
    .C(net362),
    .D(net354),
    .X(_02432_));
 sky130_fd_sc_hd__a22oi_2 _08436_ (.A1(net161),
    .A2(net362),
    .B1(net354),
    .B2(net170),
    .Y(_02433_));
 sky130_fd_sc_hd__or3_1 _08437_ (.A(_02431_),
    .B(_02432_),
    .C(_02433_),
    .X(_02434_));
 sky130_fd_sc_hd__o21ai_1 _08438_ (.A1(_02432_),
    .A2(_02433_),
    .B1(_02431_),
    .Y(_02436_));
 sky130_fd_sc_hd__o21bai_1 _08439_ (.A1(_02265_),
    .A2(_02267_),
    .B1_N(_02266_),
    .Y(_02437_));
 sky130_fd_sc_hd__and3_1 _08440_ (.A(_02434_),
    .B(_02436_),
    .C(_02437_),
    .X(_02438_));
 sky130_fd_sc_hd__a21o_1 _08441_ (.A1(_02434_),
    .A2(_02436_),
    .B1(_02437_),
    .X(_02439_));
 sky130_fd_sc_hd__and2b_1 _08442_ (.A_N(_02438_),
    .B(_02439_),
    .X(_02440_));
 sky130_fd_sc_hd__xnor2_1 _08443_ (.A(_02430_),
    .B(_02440_),
    .Y(_02441_));
 sky130_fd_sc_hd__nand2_1 _08444_ (.A(_02278_),
    .B(_02281_),
    .Y(_02442_));
 sky130_fd_sc_hd__a31o_1 _08445_ (.A1(net399),
    .A2(net595),
    .A3(_02301_),
    .B1(_02300_),
    .X(_02443_));
 sky130_fd_sc_hd__nand4_1 _08446_ (.A(net391),
    .B(net375),
    .C(net610),
    .D(net594),
    .Y(_02444_));
 sky130_fd_sc_hd__a22o_1 _08447_ (.A1(net375),
    .A2(net610),
    .B1(net594),
    .B2(net391),
    .X(_02445_));
 sky130_fd_sc_hd__a22o_1 _08448_ (.A1(net368),
    .A2(net618),
    .B1(_02444_),
    .B2(_02445_),
    .X(_02447_));
 sky130_fd_sc_hd__nand4_1 _08449_ (.A(net368),
    .B(net618),
    .C(_02444_),
    .D(_02445_),
    .Y(_02448_));
 sky130_fd_sc_hd__nand3_1 _08450_ (.A(_02443_),
    .B(_02447_),
    .C(_02448_),
    .Y(_02449_));
 sky130_fd_sc_hd__a21o_1 _08451_ (.A1(_02447_),
    .A2(_02448_),
    .B1(_02443_),
    .X(_02450_));
 sky130_fd_sc_hd__nand3_1 _08452_ (.A(_02442_),
    .B(_02449_),
    .C(_02450_),
    .Y(_02451_));
 sky130_fd_sc_hd__a21o_1 _08453_ (.A1(_02449_),
    .A2(_02450_),
    .B1(_02442_),
    .X(_02452_));
 sky130_fd_sc_hd__a21bo_1 _08454_ (.A1(_02276_),
    .A2(_02284_),
    .B1_N(_02283_),
    .X(_02453_));
 sky130_fd_sc_hd__and3_1 _08455_ (.A(_02451_),
    .B(_02452_),
    .C(_02453_),
    .X(_02454_));
 sky130_fd_sc_hd__inv_2 _08456_ (.A(_02454_),
    .Y(_02455_));
 sky130_fd_sc_hd__a21oi_1 _08457_ (.A1(_02451_),
    .A2(_02452_),
    .B1(_02453_),
    .Y(_02456_));
 sky130_fd_sc_hd__nor3_1 _08458_ (.A(_02441_),
    .B(_02454_),
    .C(_02456_),
    .Y(_02458_));
 sky130_fd_sc_hd__or3_1 _08459_ (.A(_02441_),
    .B(_02454_),
    .C(_02456_),
    .X(_02459_));
 sky130_fd_sc_hd__o21a_1 _08460_ (.A1(_02454_),
    .A2(_02456_),
    .B1(_02441_),
    .X(_02460_));
 sky130_fd_sc_hd__a211oi_1 _08461_ (.A1(_02316_),
    .A2(_02318_),
    .B1(_02458_),
    .C1(_02460_),
    .Y(_02461_));
 sky130_fd_sc_hd__o211a_1 _08462_ (.A1(_02458_),
    .A2(_02460_),
    .B1(_02316_),
    .C1(_02318_),
    .X(_02462_));
 sky130_fd_sc_hd__nor2_1 _08463_ (.A(_02461_),
    .B(_02462_),
    .Y(_02463_));
 sky130_fd_sc_hd__xnor2_1 _08464_ (.A(_02425_),
    .B(_02463_),
    .Y(_02464_));
 sky130_fd_sc_hd__nand2_1 _08465_ (.A(_02311_),
    .B(_02313_),
    .Y(_02465_));
 sky130_fd_sc_hd__a21bo_1 _08466_ (.A1(_02321_),
    .A2(_02330_),
    .B1_N(_02329_),
    .X(_02466_));
 sky130_fd_sc_hd__nand2_1 _08467_ (.A(net399),
    .B(net587),
    .Y(_02467_));
 sky130_fd_sc_hd__and4_1 _08468_ (.A(net414),
    .B(net406),
    .C(net579),
    .D(net573),
    .X(_02469_));
 sky130_fd_sc_hd__a22o_1 _08469_ (.A1(net406),
    .A2(net579),
    .B1(net573),
    .B2(net414),
    .X(_02470_));
 sky130_fd_sc_hd__and2b_1 _08470_ (.A_N(_02469_),
    .B(_02470_),
    .X(_02471_));
 sky130_fd_sc_hd__xnor2_1 _08471_ (.A(_02467_),
    .B(_02471_),
    .Y(_02472_));
 sky130_fd_sc_hd__nand2_1 _08472_ (.A(net421),
    .B(net570),
    .Y(_02473_));
 sky130_fd_sc_hd__and4_1 _08473_ (.A(net182),
    .B(net428),
    .C(net559),
    .D(net552),
    .X(_02474_));
 sky130_fd_sc_hd__a22oi_2 _08474_ (.A1(net428),
    .A2(net559),
    .B1(net552),
    .B2(net184),
    .Y(_02475_));
 sky130_fd_sc_hd__or3_1 _08475_ (.A(_02473_),
    .B(_02474_),
    .C(_02475_),
    .X(_02476_));
 sky130_fd_sc_hd__o21ai_1 _08476_ (.A1(_02474_),
    .A2(_02475_),
    .B1(_02473_),
    .Y(_02477_));
 sky130_fd_sc_hd__o21bai_1 _08477_ (.A1(_02305_),
    .A2(_02307_),
    .B1_N(_02306_),
    .Y(_02478_));
 sky130_fd_sc_hd__nand3_1 _08478_ (.A(_02476_),
    .B(_02477_),
    .C(_02478_),
    .Y(_02480_));
 sky130_fd_sc_hd__a21o_1 _08479_ (.A1(_02476_),
    .A2(_02477_),
    .B1(_02478_),
    .X(_02481_));
 sky130_fd_sc_hd__nand3_1 _08480_ (.A(_02472_),
    .B(_02480_),
    .C(_02481_),
    .Y(_02482_));
 sky130_fd_sc_hd__a21o_1 _08481_ (.A1(_02480_),
    .A2(_02481_),
    .B1(_02472_),
    .X(_02483_));
 sky130_fd_sc_hd__nand3_2 _08482_ (.A(_02466_),
    .B(_02482_),
    .C(_02483_),
    .Y(_02484_));
 sky130_fd_sc_hd__a21o_1 _08483_ (.A1(_02482_),
    .A2(_02483_),
    .B1(_02466_),
    .X(_02485_));
 sky130_fd_sc_hd__nand3_2 _08484_ (.A(_02465_),
    .B(_02484_),
    .C(_02485_),
    .Y(_02486_));
 sky130_fd_sc_hd__a21o_1 _08485_ (.A1(_02484_),
    .A2(_02485_),
    .B1(_02465_),
    .X(_02487_));
 sky130_fd_sc_hd__a22oi_1 _08486_ (.A1(net216),
    .A2(net510),
    .B1(net502),
    .B2(net229),
    .Y(_02488_));
 sky130_fd_sc_hd__and4_1 _08487_ (.A(net229),
    .B(net216),
    .C(net510),
    .D(net502),
    .X(_02489_));
 sky130_fd_sc_hd__nor2_1 _08488_ (.A(_02488_),
    .B(_02489_),
    .Y(_02491_));
 sky130_fd_sc_hd__nand2_1 _08489_ (.A(_02324_),
    .B(_02327_),
    .Y(_02492_));
 sky130_fd_sc_hd__a31o_1 _08490_ (.A1(net216),
    .A2(net524),
    .A3(_02336_),
    .B1(_02335_),
    .X(_02493_));
 sky130_fd_sc_hd__a22o_1 _08491_ (.A1(net200),
    .A2(net533),
    .B1(net523),
    .B2(net211),
    .X(_02494_));
 sky130_fd_sc_hd__nand4_1 _08492_ (.A(net211),
    .B(net200),
    .C(net533),
    .D(net523),
    .Y(_02495_));
 sky130_fd_sc_hd__a22o_1 _08493_ (.A1(net192),
    .A2(net542),
    .B1(_02494_),
    .B2(_02495_),
    .X(_02496_));
 sky130_fd_sc_hd__nand4_1 _08494_ (.A(net192),
    .B(net542),
    .C(_02494_),
    .D(_02495_),
    .Y(_02497_));
 sky130_fd_sc_hd__nand3_1 _08495_ (.A(_02493_),
    .B(_02496_),
    .C(_02497_),
    .Y(_02498_));
 sky130_fd_sc_hd__a21o_1 _08496_ (.A1(_02496_),
    .A2(_02497_),
    .B1(_02493_),
    .X(_02499_));
 sky130_fd_sc_hd__nand3_1 _08497_ (.A(_02492_),
    .B(_02498_),
    .C(_02499_),
    .Y(_02500_));
 sky130_fd_sc_hd__a21o_1 _08498_ (.A1(_02498_),
    .A2(_02499_),
    .B1(_02492_),
    .X(_02502_));
 sky130_fd_sc_hd__nand3_1 _08499_ (.A(_02491_),
    .B(_02500_),
    .C(_02502_),
    .Y(_02503_));
 sky130_fd_sc_hd__a21o_1 _08500_ (.A1(_02500_),
    .A2(_02502_),
    .B1(_02491_),
    .X(_02504_));
 sky130_fd_sc_hd__a31o_1 _08501_ (.A1(_02331_),
    .A2(_02332_),
    .A3(_02341_),
    .B1(_02340_),
    .X(_02505_));
 sky130_fd_sc_hd__and3_1 _08502_ (.A(_02503_),
    .B(_02504_),
    .C(_02505_),
    .X(_02506_));
 sky130_fd_sc_hd__nand3_1 _08503_ (.A(_02503_),
    .B(_02504_),
    .C(_02505_),
    .Y(_02507_));
 sky130_fd_sc_hd__a21o_1 _08504_ (.A1(_02503_),
    .A2(_02504_),
    .B1(_02505_),
    .X(_02508_));
 sky130_fd_sc_hd__and4_1 _08505_ (.A(_02486_),
    .B(_02487_),
    .C(_02507_),
    .D(_02508_),
    .X(_02509_));
 sky130_fd_sc_hd__a22o_1 _08506_ (.A1(_02486_),
    .A2(_02487_),
    .B1(_02507_),
    .B2(_02508_),
    .X(_02510_));
 sky130_fd_sc_hd__and2b_1 _08507_ (.A_N(_02509_),
    .B(_02510_),
    .X(_02511_));
 sky130_fd_sc_hd__a21oi_1 _08508_ (.A1(_02320_),
    .A2(_02346_),
    .B1(_02345_),
    .Y(_02513_));
 sky130_fd_sc_hd__and2b_1 _08509_ (.A_N(_02513_),
    .B(_02511_),
    .X(_02514_));
 sky130_fd_sc_hd__xnor2_1 _08510_ (.A(_02511_),
    .B(_02513_),
    .Y(_02515_));
 sky130_fd_sc_hd__xor2_1 _08511_ (.A(_02464_),
    .B(_02515_),
    .X(_02516_));
 sky130_fd_sc_hd__a21oi_1 _08512_ (.A1(_02296_),
    .A2(_02351_),
    .B1(_02350_),
    .Y(_02517_));
 sky130_fd_sc_hd__and2b_1 _08513_ (.A_N(_02517_),
    .B(_02516_),
    .X(_02518_));
 sky130_fd_sc_hd__xnor2_1 _08514_ (.A(_02516_),
    .B(_02517_),
    .Y(_02519_));
 sky130_fd_sc_hd__xnor2_1 _08515_ (.A(_02423_),
    .B(_02519_),
    .Y(_02520_));
 sky130_fd_sc_hd__a21oi_1 _08516_ (.A1(_02257_),
    .A2(_02355_),
    .B1(_02354_),
    .Y(_02521_));
 sky130_fd_sc_hd__or2_1 _08517_ (.A(_02520_),
    .B(_02521_),
    .X(_02522_));
 sky130_fd_sc_hd__xnor2_1 _08518_ (.A(_02520_),
    .B(_02521_),
    .Y(_02524_));
 sky130_fd_sc_hd__xnor2_1 _08519_ (.A(_02377_),
    .B(_02524_),
    .Y(_02525_));
 sky130_fd_sc_hd__a21oi_1 _08520_ (.A1(_02212_),
    .A2(_02360_),
    .B1(_02358_),
    .Y(_02526_));
 sky130_fd_sc_hd__and2b_1 _08521_ (.A_N(_02526_),
    .B(_02525_),
    .X(_02527_));
 sky130_fd_sc_hd__xnor2_1 _08522_ (.A(_02525_),
    .B(_02526_),
    .Y(_02528_));
 sky130_fd_sc_hd__xnor2_1 _08523_ (.A(_02376_),
    .B(_02528_),
    .Y(_02529_));
 sky130_fd_sc_hd__a21o_1 _08524_ (.A1(_02364_),
    .A2(_02366_),
    .B1(_02529_),
    .X(_02530_));
 sky130_fd_sc_hd__inv_2 _08525_ (.A(_02530_),
    .Y(_02531_));
 sky130_fd_sc_hd__and3_1 _08526_ (.A(_02364_),
    .B(_02366_),
    .C(_02529_),
    .X(_02532_));
 sky130_fd_sc_hd__nor2_1 _08527_ (.A(_02531_),
    .B(_02532_),
    .Y(_02533_));
 sky130_fd_sc_hd__a21bo_1 _08528_ (.A1(_02371_),
    .A2(_02375_),
    .B1_N(_02369_),
    .X(_02535_));
 sky130_fd_sc_hd__xor2_1 _08529_ (.A(_02533_),
    .B(_02535_),
    .X(net93));
 sky130_fd_sc_hd__a31o_1 _08530_ (.A1(net488),
    .A2(net247),
    .A3(_02396_),
    .B1(_02395_),
    .X(_02536_));
 sky130_fd_sc_hd__o21ai_1 _08531_ (.A1(_02379_),
    .A2(_02422_),
    .B1(_02421_),
    .Y(_02537_));
 sky130_fd_sc_hd__a21bo_1 _08532_ (.A1(_02398_),
    .A2(_02418_),
    .B1_N(_02417_),
    .X(_02538_));
 sky130_fd_sc_hd__o21bai_1 _08533_ (.A1(_02425_),
    .A2(_02462_),
    .B1_N(_02461_),
    .Y(_02539_));
 sky130_fd_sc_hd__and4_1 _08534_ (.A(net449),
    .B(net442),
    .C(net280),
    .D(net273),
    .X(_02540_));
 sky130_fd_sc_hd__a22oi_1 _08535_ (.A1(net442),
    .A2(net280),
    .B1(net273),
    .B2(net449),
    .Y(_02541_));
 sky130_fd_sc_hd__o2bb2a_1 _08536_ (.A1_N(net459),
    .A2_N(net263),
    .B1(_02540_),
    .B2(_02541_),
    .X(_02542_));
 sky130_fd_sc_hd__and4bb_1 _08537_ (.A_N(_02540_),
    .B_N(_02541_),
    .C(net459),
    .D(net264),
    .X(_02543_));
 sky130_fd_sc_hd__nor2_1 _08538_ (.A(_02542_),
    .B(_02543_),
    .Y(_02545_));
 sky130_fd_sc_hd__nor2_1 _08539_ (.A(_02382_),
    .B(_02385_),
    .Y(_02546_));
 sky130_fd_sc_hd__and2b_1 _08540_ (.A_N(_02546_),
    .B(_02545_),
    .X(_02547_));
 sky130_fd_sc_hd__xnor2_1 _08541_ (.A(_02545_),
    .B(_02546_),
    .Y(_02548_));
 sky130_fd_sc_hd__and2_1 _08542_ (.A(net473),
    .B(net252),
    .X(_02549_));
 sky130_fd_sc_hd__xnor2_1 _08543_ (.A(_02548_),
    .B(_02549_),
    .Y(_02550_));
 sky130_fd_sc_hd__and3_1 _08544_ (.A(_02388_),
    .B(_02392_),
    .C(_02550_),
    .X(_02551_));
 sky130_fd_sc_hd__a21oi_1 _08545_ (.A1(_02388_),
    .A2(_02392_),
    .B1(_02550_),
    .Y(_02552_));
 sky130_fd_sc_hd__nor2_1 _08546_ (.A(_02551_),
    .B(_02552_),
    .Y(_02553_));
 sky130_fd_sc_hd__nand2_1 _08547_ (.A(net481),
    .B(net247),
    .Y(_02554_));
 sky130_fd_sc_hd__xnor2_1 _08548_ (.A(_02553_),
    .B(_02554_),
    .Y(_02556_));
 sky130_fd_sc_hd__a21o_1 _08549_ (.A1(_02430_),
    .A2(_02439_),
    .B1(_02438_),
    .X(_02557_));
 sky130_fd_sc_hd__nand2_1 _08550_ (.A(_02403_),
    .B(_02406_),
    .Y(_02558_));
 sky130_fd_sc_hd__a31o_1 _08551_ (.A1(net382),
    .A2(net316),
    .A3(_02427_),
    .B1(_02426_),
    .X(_02559_));
 sky130_fd_sc_hd__nand4_2 _08552_ (.A(net463),
    .B(net382),
    .C(net308),
    .D(net294),
    .Y(_02560_));
 sky130_fd_sc_hd__a22o_1 _08553_ (.A1(net382),
    .A2(net308),
    .B1(net294),
    .B2(net463),
    .X(_02561_));
 sky130_fd_sc_hd__a22o_1 _08554_ (.A1(net543),
    .A2(net287),
    .B1(_02560_),
    .B2(_02561_),
    .X(_02562_));
 sky130_fd_sc_hd__nand4_2 _08555_ (.A(net543),
    .B(net287),
    .C(_02560_),
    .D(_02561_),
    .Y(_02563_));
 sky130_fd_sc_hd__nand3_2 _08556_ (.A(_02559_),
    .B(_02562_),
    .C(_02563_),
    .Y(_02564_));
 sky130_fd_sc_hd__a21o_1 _08557_ (.A1(_02562_),
    .A2(_02563_),
    .B1(_02559_),
    .X(_02565_));
 sky130_fd_sc_hd__nand3_2 _08558_ (.A(_02558_),
    .B(_02564_),
    .C(_02565_),
    .Y(_02567_));
 sky130_fd_sc_hd__a21o_1 _08559_ (.A1(_02564_),
    .A2(_02565_),
    .B1(_02558_),
    .X(_02568_));
 sky130_fd_sc_hd__and3_1 _08560_ (.A(_02557_),
    .B(_02567_),
    .C(_02568_),
    .X(_02569_));
 sky130_fd_sc_hd__a21oi_1 _08561_ (.A1(_02567_),
    .A2(_02568_),
    .B1(_02557_),
    .Y(_02570_));
 sky130_fd_sc_hd__a211oi_1 _08562_ (.A1(_02407_),
    .A2(_02409_),
    .B1(_02569_),
    .C1(_02570_),
    .Y(_02571_));
 sky130_fd_sc_hd__a211o_1 _08563_ (.A1(_02407_),
    .A2(_02409_),
    .B1(_02569_),
    .C1(_02570_),
    .X(_02572_));
 sky130_fd_sc_hd__o211ai_1 _08564_ (.A1(_02569_),
    .A2(_02570_),
    .B1(_02407_),
    .C1(_02409_),
    .Y(_02573_));
 sky130_fd_sc_hd__o211a_1 _08565_ (.A1(_02411_),
    .A2(_02414_),
    .B1(_02572_),
    .C1(_02573_),
    .X(_02574_));
 sky130_fd_sc_hd__a211oi_1 _08566_ (.A1(_02572_),
    .A2(_02573_),
    .B1(_02411_),
    .C1(_02414_),
    .Y(_02575_));
 sky130_fd_sc_hd__nor2_1 _08567_ (.A(_02574_),
    .B(_02575_),
    .Y(_02576_));
 sky130_fd_sc_hd__and2_1 _08568_ (.A(_02556_),
    .B(_02576_),
    .X(_02578_));
 sky130_fd_sc_hd__xnor2_1 _08569_ (.A(_02556_),
    .B(_02576_),
    .Y(_02579_));
 sky130_fd_sc_hd__and2b_1 _08570_ (.A_N(_02579_),
    .B(_02539_),
    .X(_02580_));
 sky130_fd_sc_hd__xnor2_1 _08571_ (.A(_02539_),
    .B(_02579_),
    .Y(_02581_));
 sky130_fd_sc_hd__xor2_1 _08572_ (.A(_02538_),
    .B(_02581_),
    .X(_02582_));
 sky130_fd_sc_hd__and4_1 _08573_ (.A(net221),
    .B(net177),
    .C(net330),
    .D(net323),
    .X(_02583_));
 sky130_fd_sc_hd__a22o_1 _08574_ (.A1(net177),
    .A2(net330),
    .B1(net323),
    .B2(net221),
    .X(_02584_));
 sky130_fd_sc_hd__and2b_1 _08575_ (.A_N(_02583_),
    .B(_02584_),
    .X(_02585_));
 sky130_fd_sc_hd__nand2_1 _08576_ (.A(net298),
    .B(net316),
    .Y(_02586_));
 sky130_fd_sc_hd__xnor2_1 _08577_ (.A(_02585_),
    .B(_02586_),
    .Y(_02587_));
 sky130_fd_sc_hd__nand4_1 _08578_ (.A(net161),
    .B(net619),
    .C(net362),
    .D(net354),
    .Y(_02589_));
 sky130_fd_sc_hd__a22o_1 _08579_ (.A1(net619),
    .A2(net362),
    .B1(net354),
    .B2(net161),
    .X(_02590_));
 sky130_fd_sc_hd__and2_1 _08580_ (.A(net169),
    .B(net339),
    .X(_02591_));
 sky130_fd_sc_hd__a21o_1 _08581_ (.A1(_02589_),
    .A2(_02590_),
    .B1(_02591_),
    .X(_02592_));
 sky130_fd_sc_hd__nand3_1 _08582_ (.A(_02589_),
    .B(_02590_),
    .C(_02591_),
    .Y(_02593_));
 sky130_fd_sc_hd__o21bai_1 _08583_ (.A1(_02431_),
    .A2(_02433_),
    .B1_N(_02432_),
    .Y(_02594_));
 sky130_fd_sc_hd__and3_1 _08584_ (.A(_02592_),
    .B(_02593_),
    .C(_02594_),
    .X(_02595_));
 sky130_fd_sc_hd__a21o_1 _08585_ (.A1(_02592_),
    .A2(_02593_),
    .B1(_02594_),
    .X(_02596_));
 sky130_fd_sc_hd__and2b_1 _08586_ (.A_N(_02595_),
    .B(_02596_),
    .X(_02597_));
 sky130_fd_sc_hd__xnor2_1 _08587_ (.A(_02587_),
    .B(_02597_),
    .Y(_02598_));
 sky130_fd_sc_hd__nand2_1 _08588_ (.A(_02444_),
    .B(_02448_),
    .Y(_02600_));
 sky130_fd_sc_hd__a31o_1 _08589_ (.A1(net399),
    .A2(net587),
    .A3(_02470_),
    .B1(_02469_),
    .X(_02601_));
 sky130_fd_sc_hd__nand4_1 _08590_ (.A(net391),
    .B(net375),
    .C(net595),
    .D(net587),
    .Y(_02602_));
 sky130_fd_sc_hd__a22o_1 _08591_ (.A1(net375),
    .A2(net594),
    .B1(net587),
    .B2(net391),
    .X(_02603_));
 sky130_fd_sc_hd__a22o_1 _08592_ (.A1(net368),
    .A2(net611),
    .B1(_02602_),
    .B2(_02603_),
    .X(_02604_));
 sky130_fd_sc_hd__nand4_1 _08593_ (.A(net368),
    .B(net611),
    .C(_02602_),
    .D(_02603_),
    .Y(_02605_));
 sky130_fd_sc_hd__nand3_1 _08594_ (.A(_02601_),
    .B(_02604_),
    .C(_02605_),
    .Y(_02606_));
 sky130_fd_sc_hd__a21o_1 _08595_ (.A1(_02604_),
    .A2(_02605_),
    .B1(_02601_),
    .X(_02607_));
 sky130_fd_sc_hd__nand3_1 _08596_ (.A(_02600_),
    .B(_02606_),
    .C(_02607_),
    .Y(_02608_));
 sky130_fd_sc_hd__a21o_1 _08597_ (.A1(_02606_),
    .A2(_02607_),
    .B1(_02600_),
    .X(_02609_));
 sky130_fd_sc_hd__a21bo_1 _08598_ (.A1(_02442_),
    .A2(_02450_),
    .B1_N(_02449_),
    .X(_02611_));
 sky130_fd_sc_hd__and3_1 _08599_ (.A(_02608_),
    .B(_02609_),
    .C(_02611_),
    .X(_02612_));
 sky130_fd_sc_hd__inv_2 _08600_ (.A(_02612_),
    .Y(_02613_));
 sky130_fd_sc_hd__a21oi_1 _08601_ (.A1(_02608_),
    .A2(_02609_),
    .B1(_02611_),
    .Y(_02614_));
 sky130_fd_sc_hd__nor3_1 _08602_ (.A(_02598_),
    .B(_02612_),
    .C(_02614_),
    .Y(_02615_));
 sky130_fd_sc_hd__or3_2 _08603_ (.A(_02598_),
    .B(_02612_),
    .C(_02614_),
    .X(_02616_));
 sky130_fd_sc_hd__o21a_1 _08604_ (.A1(_02612_),
    .A2(_02614_),
    .B1(_02598_),
    .X(_02617_));
 sky130_fd_sc_hd__a211oi_4 _08605_ (.A1(_02484_),
    .A2(_02486_),
    .B1(net157),
    .C1(_02617_),
    .Y(_02618_));
 sky130_fd_sc_hd__o211a_1 _08606_ (.A1(_02615_),
    .A2(_02617_),
    .B1(_02484_),
    .C1(_02486_),
    .X(_02619_));
 sky130_fd_sc_hd__a211oi_2 _08607_ (.A1(_02455_),
    .A2(_02459_),
    .B1(_02618_),
    .C1(_02619_),
    .Y(_02620_));
 sky130_fd_sc_hd__o211a_1 _08608_ (.A1(_02618_),
    .A2(_02619_),
    .B1(_02455_),
    .C1(_02459_),
    .X(_02622_));
 sky130_fd_sc_hd__nand2_1 _08609_ (.A(_02480_),
    .B(_02482_),
    .Y(_02623_));
 sky130_fd_sc_hd__a21bo_1 _08610_ (.A1(_02492_),
    .A2(_02499_),
    .B1_N(_02498_),
    .X(_02624_));
 sky130_fd_sc_hd__and4_1 _08611_ (.A(net414),
    .B(net406),
    .C(net573),
    .D(net566),
    .X(_02625_));
 sky130_fd_sc_hd__a22o_1 _08612_ (.A1(net406),
    .A2(net573),
    .B1(net566),
    .B2(net414),
    .X(_02626_));
 sky130_fd_sc_hd__and2b_1 _08613_ (.A_N(_02625_),
    .B(_02626_),
    .X(_02627_));
 sky130_fd_sc_hd__nand2_1 _08614_ (.A(net399),
    .B(net579),
    .Y(_02628_));
 sky130_fd_sc_hd__xnor2_1 _08615_ (.A(_02627_),
    .B(_02628_),
    .Y(_02629_));
 sky130_fd_sc_hd__nand4_1 _08616_ (.A(net184),
    .B(net428),
    .C(net552),
    .D(net538),
    .Y(_02630_));
 sky130_fd_sc_hd__a22o_1 _08617_ (.A1(net428),
    .A2(net553),
    .B1(net538),
    .B2(net184),
    .X(_02631_));
 sky130_fd_sc_hd__and2_1 _08618_ (.A(net421),
    .B(net563),
    .X(_02633_));
 sky130_fd_sc_hd__a21o_1 _08619_ (.A1(_02630_),
    .A2(_02631_),
    .B1(_02633_),
    .X(_02634_));
 sky130_fd_sc_hd__nand3_1 _08620_ (.A(_02630_),
    .B(_02631_),
    .C(_02633_),
    .Y(_02635_));
 sky130_fd_sc_hd__o21bai_1 _08621_ (.A1(_02473_),
    .A2(_02475_),
    .B1_N(_02474_),
    .Y(_02636_));
 sky130_fd_sc_hd__nand3_1 _08622_ (.A(_02634_),
    .B(_02635_),
    .C(_02636_),
    .Y(_02637_));
 sky130_fd_sc_hd__a21o_1 _08623_ (.A1(_02634_),
    .A2(_02635_),
    .B1(_02636_),
    .X(_02638_));
 sky130_fd_sc_hd__nand3_1 _08624_ (.A(_02629_),
    .B(_02637_),
    .C(_02638_),
    .Y(_02639_));
 sky130_fd_sc_hd__a21o_1 _08625_ (.A1(_02637_),
    .A2(_02638_),
    .B1(_02629_),
    .X(_02640_));
 sky130_fd_sc_hd__nand3_2 _08626_ (.A(_02624_),
    .B(_02639_),
    .C(_02640_),
    .Y(_02641_));
 sky130_fd_sc_hd__a21o_1 _08627_ (.A1(_02639_),
    .A2(_02640_),
    .B1(_02624_),
    .X(_02642_));
 sky130_fd_sc_hd__nand3_2 _08628_ (.A(_02623_),
    .B(_02641_),
    .C(_02642_),
    .Y(_02644_));
 sky130_fd_sc_hd__a21o_1 _08629_ (.A1(_02641_),
    .A2(_02642_),
    .B1(_02623_),
    .X(_02645_));
 sky130_fd_sc_hd__nand2_1 _08630_ (.A(_02495_),
    .B(_02497_),
    .Y(_02646_));
 sky130_fd_sc_hd__and2_1 _08631_ (.A(net200),
    .B(net510),
    .X(_02647_));
 sky130_fd_sc_hd__nand2_1 _08632_ (.A(net206),
    .B(net510),
    .Y(_02648_));
 sky130_fd_sc_hd__nand4_1 _08633_ (.A(net211),
    .B(net200),
    .C(net523),
    .D(net509),
    .Y(_02649_));
 sky130_fd_sc_hd__a22o_1 _08634_ (.A1(net202),
    .A2(net523),
    .B1(net510),
    .B2(net211),
    .X(_02650_));
 sky130_fd_sc_hd__nand2_1 _08635_ (.A(net192),
    .B(net533),
    .Y(_02651_));
 sky130_fd_sc_hd__a21bo_1 _08636_ (.A1(_02649_),
    .A2(_02650_),
    .B1_N(_02651_),
    .X(_02652_));
 sky130_fd_sc_hd__nand3b_1 _08637_ (.A_N(_02651_),
    .B(_02650_),
    .C(_02649_),
    .Y(_02653_));
 sky130_fd_sc_hd__nand3_1 _08638_ (.A(_02489_),
    .B(_02652_),
    .C(_02653_),
    .Y(_02655_));
 sky130_fd_sc_hd__a21o_1 _08639_ (.A1(_02652_),
    .A2(_02653_),
    .B1(_02489_),
    .X(_02656_));
 sky130_fd_sc_hd__nand3_1 _08640_ (.A(_02646_),
    .B(_02655_),
    .C(_02656_),
    .Y(_02657_));
 sky130_fd_sc_hd__a21o_1 _08641_ (.A1(_02655_),
    .A2(_02656_),
    .B1(_02646_),
    .X(_02658_));
 sky130_fd_sc_hd__nand4_2 _08642_ (.A(net218),
    .B(net502),
    .C(_02657_),
    .D(_02658_),
    .Y(_02659_));
 sky130_fd_sc_hd__a22o_1 _08643_ (.A1(net218),
    .A2(net502),
    .B1(_02657_),
    .B2(_02658_),
    .X(_02660_));
 sky130_fd_sc_hd__nand3b_2 _08644_ (.A_N(_02503_),
    .B(_02659_),
    .C(_02660_),
    .Y(_02661_));
 sky130_fd_sc_hd__a21bo_1 _08645_ (.A1(_02659_),
    .A2(_02660_),
    .B1_N(_02503_),
    .X(_02662_));
 sky130_fd_sc_hd__nand4_2 _08646_ (.A(_02644_),
    .B(_02645_),
    .C(_02661_),
    .D(_02662_),
    .Y(_02663_));
 sky130_fd_sc_hd__a22o_1 _08647_ (.A1(_02644_),
    .A2(_02645_),
    .B1(_02661_),
    .B2(_02662_),
    .X(_02664_));
 sky130_fd_sc_hd__o211a_1 _08648_ (.A1(_02506_),
    .A2(_02509_),
    .B1(_02663_),
    .C1(_02664_),
    .X(_02666_));
 sky130_fd_sc_hd__a211oi_1 _08649_ (.A1(_02663_),
    .A2(_02664_),
    .B1(_02506_),
    .C1(_02509_),
    .Y(_02667_));
 sky130_fd_sc_hd__nor4_1 _08650_ (.A(_02620_),
    .B(_02622_),
    .C(_02666_),
    .D(_02667_),
    .Y(_02668_));
 sky130_fd_sc_hd__o22a_1 _08651_ (.A1(_02620_),
    .A2(_02622_),
    .B1(_02666_),
    .B2(_02667_),
    .X(_02669_));
 sky130_fd_sc_hd__nor2_1 _08652_ (.A(_02668_),
    .B(_02669_),
    .Y(_02670_));
 sky130_fd_sc_hd__a21o_1 _08653_ (.A1(_02464_),
    .A2(_02515_),
    .B1(_02514_),
    .X(_02671_));
 sky130_fd_sc_hd__nand2_1 _08654_ (.A(_02670_),
    .B(_02671_),
    .Y(_02672_));
 sky130_fd_sc_hd__xor2_1 _08655_ (.A(_02670_),
    .B(_02671_),
    .X(_02673_));
 sky130_fd_sc_hd__xnor2_1 _08656_ (.A(_02582_),
    .B(_02673_),
    .Y(_02674_));
 sky130_fd_sc_hd__a21oi_1 _08657_ (.A1(_02423_),
    .A2(_02519_),
    .B1(_02518_),
    .Y(_02675_));
 sky130_fd_sc_hd__nor2_1 _08658_ (.A(_02674_),
    .B(_02675_),
    .Y(_02677_));
 sky130_fd_sc_hd__nand2_1 _08659_ (.A(_02674_),
    .B(_02675_),
    .Y(_02678_));
 sky130_fd_sc_hd__xnor2_1 _08660_ (.A(_02674_),
    .B(_02675_),
    .Y(_02679_));
 sky130_fd_sc_hd__xnor2_1 _08661_ (.A(_02537_),
    .B(_02679_),
    .Y(_02680_));
 sky130_fd_sc_hd__o21ai_1 _08662_ (.A1(_02378_),
    .A2(_02524_),
    .B1(_02522_),
    .Y(_02681_));
 sky130_fd_sc_hd__nand2_1 _08663_ (.A(_02680_),
    .B(_02681_),
    .Y(_02682_));
 sky130_fd_sc_hd__xor2_1 _08664_ (.A(_02680_),
    .B(_02681_),
    .X(_02683_));
 sky130_fd_sc_hd__nand2_1 _08665_ (.A(_02536_),
    .B(_02683_),
    .Y(_02684_));
 sky130_fd_sc_hd__xnor2_1 _08666_ (.A(_02536_),
    .B(_02683_),
    .Y(_02685_));
 sky130_fd_sc_hd__a21oi_1 _08667_ (.A1(_02376_),
    .A2(_02528_),
    .B1(_02527_),
    .Y(_02686_));
 sky130_fd_sc_hd__or2_1 _08668_ (.A(_02685_),
    .B(_02686_),
    .X(_02688_));
 sky130_fd_sc_hd__xor2_1 _08669_ (.A(_02685_),
    .B(_02686_),
    .X(_02689_));
 sky130_fd_sc_hd__or3b_1 _08670_ (.A(_02532_),
    .B(_02372_),
    .C_N(_02530_),
    .X(_02690_));
 sky130_fd_sc_hd__o221a_1 _08671_ (.A1(_02369_),
    .A2(_02532_),
    .B1(_02690_),
    .B2(_02373_),
    .C1(_02530_),
    .X(_02691_));
 sky130_fd_sc_hd__or4b_2 _08672_ (.A(_02207_),
    .B(_02208_),
    .C(_02690_),
    .D_N(_02035_),
    .X(_02692_));
 sky130_fd_sc_hd__o21ai_2 _08673_ (.A1(_02046_),
    .A2(_02692_),
    .B1(_02691_),
    .Y(_02693_));
 sky130_fd_sc_hd__xor2_1 _08674_ (.A(_02689_),
    .B(_02693_),
    .X(net94));
 sky130_fd_sc_hd__a31o_1 _08675_ (.A1(net481),
    .A2(net247),
    .A3(_02553_),
    .B1(_02552_),
    .X(_02694_));
 sky130_fd_sc_hd__a21o_1 _08676_ (.A1(_02538_),
    .A2(_02581_),
    .B1(_02580_),
    .X(_02695_));
 sky130_fd_sc_hd__and4_1 _08677_ (.A(net543),
    .B(net442),
    .C(net281),
    .D(net272),
    .X(_02696_));
 sky130_fd_sc_hd__a22oi_1 _08678_ (.A1(net543),
    .A2(net281),
    .B1(net272),
    .B2(net442),
    .Y(_02698_));
 sky130_fd_sc_hd__o2bb2a_1 _08679_ (.A1_N(net449),
    .A2_N(net263),
    .B1(_02696_),
    .B2(_02698_),
    .X(_02699_));
 sky130_fd_sc_hd__and4bb_1 _08680_ (.A_N(_02696_),
    .B_N(_02698_),
    .C(net449),
    .D(net263),
    .X(_02700_));
 sky130_fd_sc_hd__nor2_1 _08681_ (.A(_02699_),
    .B(_02700_),
    .Y(_02701_));
 sky130_fd_sc_hd__nor2_1 _08682_ (.A(_02540_),
    .B(_02543_),
    .Y(_02702_));
 sky130_fd_sc_hd__and2b_1 _08683_ (.A_N(_02702_),
    .B(_02701_),
    .X(_02703_));
 sky130_fd_sc_hd__xnor2_1 _08684_ (.A(_02701_),
    .B(_02702_),
    .Y(_02704_));
 sky130_fd_sc_hd__and2_1 _08685_ (.A(net459),
    .B(net253),
    .X(_02705_));
 sky130_fd_sc_hd__xnor2_1 _08686_ (.A(_02704_),
    .B(_02705_),
    .Y(_02706_));
 sky130_fd_sc_hd__a21oi_1 _08687_ (.A1(_02548_),
    .A2(_02549_),
    .B1(_02547_),
    .Y(_02707_));
 sky130_fd_sc_hd__xnor2_1 _08688_ (.A(_02706_),
    .B(_02707_),
    .Y(_02709_));
 sky130_fd_sc_hd__nand2_1 _08689_ (.A(net477),
    .B(net248),
    .Y(_02710_));
 sky130_fd_sc_hd__or2_1 _08690_ (.A(_02709_),
    .B(_02710_),
    .X(_02711_));
 sky130_fd_sc_hd__xor2_1 _08691_ (.A(_02709_),
    .B(_02710_),
    .X(_02712_));
 sky130_fd_sc_hd__a21o_1 _08692_ (.A1(_02587_),
    .A2(_02596_),
    .B1(_02595_),
    .X(_02713_));
 sky130_fd_sc_hd__nand2_1 _08693_ (.A(_02560_),
    .B(_02563_),
    .Y(_02714_));
 sky130_fd_sc_hd__a31o_1 _08694_ (.A1(net298),
    .A2(net316),
    .A3(_02584_),
    .B1(_02583_),
    .X(_02715_));
 sky130_fd_sc_hd__nand4_2 _08695_ (.A(net381),
    .B(net298),
    .C(net308),
    .D(net294),
    .Y(_02716_));
 sky130_fd_sc_hd__a22o_1 _08696_ (.A1(net298),
    .A2(net308),
    .B1(net294),
    .B2(net382),
    .X(_02717_));
 sky130_fd_sc_hd__a22o_1 _08697_ (.A1(net464),
    .A2(net287),
    .B1(_02716_),
    .B2(_02717_),
    .X(_02718_));
 sky130_fd_sc_hd__nand4_2 _08698_ (.A(net464),
    .B(net287),
    .C(_02716_),
    .D(_02717_),
    .Y(_02720_));
 sky130_fd_sc_hd__nand3_2 _08699_ (.A(_02715_),
    .B(_02718_),
    .C(_02720_),
    .Y(_02721_));
 sky130_fd_sc_hd__a21o_1 _08700_ (.A1(_02718_),
    .A2(_02720_),
    .B1(_02715_),
    .X(_02722_));
 sky130_fd_sc_hd__nand3_2 _08701_ (.A(_02714_),
    .B(_02721_),
    .C(_02722_),
    .Y(_02723_));
 sky130_fd_sc_hd__a21o_1 _08702_ (.A1(_02721_),
    .A2(_02722_),
    .B1(_02714_),
    .X(_02724_));
 sky130_fd_sc_hd__and3_2 _08703_ (.A(_02713_),
    .B(_02723_),
    .C(_02724_),
    .X(_02725_));
 sky130_fd_sc_hd__a21oi_2 _08704_ (.A1(_02723_),
    .A2(_02724_),
    .B1(_02713_),
    .Y(_02726_));
 sky130_fd_sc_hd__a211oi_2 _08705_ (.A1(_02564_),
    .A2(_02567_),
    .B1(_02725_),
    .C1(_02726_),
    .Y(_02727_));
 sky130_fd_sc_hd__a211o_1 _08706_ (.A1(_02564_),
    .A2(_02567_),
    .B1(_02725_),
    .C1(_02726_),
    .X(_02728_));
 sky130_fd_sc_hd__o211ai_2 _08707_ (.A1(_02725_),
    .A2(_02726_),
    .B1(_02564_),
    .C1(_02567_),
    .Y(_02729_));
 sky130_fd_sc_hd__o211ai_2 _08708_ (.A1(_02569_),
    .A2(_02571_),
    .B1(_02728_),
    .C1(_02729_),
    .Y(_02731_));
 sky130_fd_sc_hd__inv_2 _08709_ (.A(_02731_),
    .Y(_02732_));
 sky130_fd_sc_hd__a211o_1 _08710_ (.A1(_02728_),
    .A2(_02729_),
    .B1(_02569_),
    .C1(_02571_),
    .X(_02733_));
 sky130_fd_sc_hd__and3_1 _08711_ (.A(_02712_),
    .B(_02731_),
    .C(_02733_),
    .X(_02734_));
 sky130_fd_sc_hd__nand3_1 _08712_ (.A(_02712_),
    .B(_02731_),
    .C(_02733_),
    .Y(_02735_));
 sky130_fd_sc_hd__a21o_1 _08713_ (.A1(_02731_),
    .A2(_02733_),
    .B1(_02712_),
    .X(_02736_));
 sky130_fd_sc_hd__o211a_1 _08714_ (.A1(_02618_),
    .A2(_02620_),
    .B1(_02735_),
    .C1(_02736_),
    .X(_02737_));
 sky130_fd_sc_hd__o211ai_1 _08715_ (.A1(_02618_),
    .A2(_02620_),
    .B1(_02735_),
    .C1(_02736_),
    .Y(_02738_));
 sky130_fd_sc_hd__a211o_1 _08716_ (.A1(_02735_),
    .A2(_02736_),
    .B1(_02618_),
    .C1(_02620_),
    .X(_02739_));
 sky130_fd_sc_hd__o211a_1 _08717_ (.A1(_02574_),
    .A2(_02578_),
    .B1(_02738_),
    .C1(_02739_),
    .X(_02740_));
 sky130_fd_sc_hd__a211oi_1 _08718_ (.A1(_02738_),
    .A2(_02739_),
    .B1(_02574_),
    .C1(_02578_),
    .Y(_02742_));
 sky130_fd_sc_hd__and4_1 _08719_ (.A(net177),
    .B(net169),
    .C(net328),
    .D(net320),
    .X(_02743_));
 sky130_fd_sc_hd__a22o_1 _08720_ (.A1(net169),
    .A2(net328),
    .B1(net320),
    .B2(net177),
    .X(_02744_));
 sky130_fd_sc_hd__and2b_1 _08721_ (.A_N(_02743_),
    .B(_02744_),
    .X(_02745_));
 sky130_fd_sc_hd__nand2_1 _08722_ (.A(net221),
    .B(net313),
    .Y(_02746_));
 sky130_fd_sc_hd__xnor2_1 _08723_ (.A(_02745_),
    .B(_02746_),
    .Y(_02747_));
 sky130_fd_sc_hd__nand4_1 _08724_ (.A(net623),
    .B(net358),
    .C(net611),
    .D(net350),
    .Y(_02748_));
 sky130_fd_sc_hd__a22o_1 _08725_ (.A1(net358),
    .A2(net611),
    .B1(net350),
    .B2(net623),
    .X(_02749_));
 sky130_fd_sc_hd__and2_1 _08726_ (.A(net161),
    .B(net335),
    .X(_02750_));
 sky130_fd_sc_hd__a21o_1 _08727_ (.A1(_02748_),
    .A2(_02749_),
    .B1(_02750_),
    .X(_02751_));
 sky130_fd_sc_hd__nand3_1 _08728_ (.A(_02748_),
    .B(_02749_),
    .C(_02750_),
    .Y(_02753_));
 sky130_fd_sc_hd__a21bo_1 _08729_ (.A1(_02590_),
    .A2(_02591_),
    .B1_N(_02589_),
    .X(_02754_));
 sky130_fd_sc_hd__and3_1 _08730_ (.A(_02751_),
    .B(_02753_),
    .C(_02754_),
    .X(_02755_));
 sky130_fd_sc_hd__a21o_1 _08731_ (.A1(_02751_),
    .A2(_02753_),
    .B1(_02754_),
    .X(_02756_));
 sky130_fd_sc_hd__and2b_1 _08732_ (.A_N(_02755_),
    .B(_02756_),
    .X(_02757_));
 sky130_fd_sc_hd__xnor2_1 _08733_ (.A(_02747_),
    .B(_02757_),
    .Y(_02758_));
 sky130_fd_sc_hd__nand2_1 _08734_ (.A(_02602_),
    .B(_02605_),
    .Y(_02759_));
 sky130_fd_sc_hd__a31o_1 _08735_ (.A1(net399),
    .A2(net579),
    .A3(_02626_),
    .B1(_02625_),
    .X(_02760_));
 sky130_fd_sc_hd__nand4_1 _08736_ (.A(net390),
    .B(net374),
    .C(net588),
    .D(net580),
    .Y(_02761_));
 sky130_fd_sc_hd__a22o_1 _08737_ (.A1(net374),
    .A2(net588),
    .B1(net580),
    .B2(net390),
    .X(_02762_));
 sky130_fd_sc_hd__a22o_1 _08738_ (.A1(net366),
    .A2(net595),
    .B1(_02761_),
    .B2(_02762_),
    .X(_02764_));
 sky130_fd_sc_hd__nand4_1 _08739_ (.A(net366),
    .B(net595),
    .C(_02761_),
    .D(_02762_),
    .Y(_02765_));
 sky130_fd_sc_hd__nand3_1 _08740_ (.A(_02760_),
    .B(_02764_),
    .C(_02765_),
    .Y(_02766_));
 sky130_fd_sc_hd__a21o_1 _08741_ (.A1(_02764_),
    .A2(_02765_),
    .B1(_02760_),
    .X(_02767_));
 sky130_fd_sc_hd__nand3_1 _08742_ (.A(_02759_),
    .B(_02766_),
    .C(_02767_),
    .Y(_02768_));
 sky130_fd_sc_hd__a21o_1 _08743_ (.A1(_02766_),
    .A2(_02767_),
    .B1(_02759_),
    .X(_02769_));
 sky130_fd_sc_hd__a21bo_1 _08744_ (.A1(_02600_),
    .A2(_02607_),
    .B1_N(_02606_),
    .X(_02770_));
 sky130_fd_sc_hd__and3_1 _08745_ (.A(_02768_),
    .B(_02769_),
    .C(_02770_),
    .X(_02771_));
 sky130_fd_sc_hd__inv_2 _08746_ (.A(_02771_),
    .Y(_02772_));
 sky130_fd_sc_hd__a21oi_1 _08747_ (.A1(_02768_),
    .A2(_02769_),
    .B1(_02770_),
    .Y(_02773_));
 sky130_fd_sc_hd__nor3_1 _08748_ (.A(_02758_),
    .B(_02771_),
    .C(_02773_),
    .Y(_02775_));
 sky130_fd_sc_hd__or3_2 _08749_ (.A(_02758_),
    .B(_02771_),
    .C(_02773_),
    .X(_02776_));
 sky130_fd_sc_hd__o21a_1 _08750_ (.A1(_02771_),
    .A2(_02773_),
    .B1(_02758_),
    .X(_02777_));
 sky130_fd_sc_hd__a211oi_4 _08751_ (.A1(_02641_),
    .A2(_02644_),
    .B1(net156),
    .C1(_02777_),
    .Y(_02778_));
 sky130_fd_sc_hd__o211a_1 _08752_ (.A1(_02775_),
    .A2(_02777_),
    .B1(_02641_),
    .C1(_02644_),
    .X(_02779_));
 sky130_fd_sc_hd__a211oi_4 _08753_ (.A1(_02613_),
    .A2(_02616_),
    .B1(_02778_),
    .C1(_02779_),
    .Y(_02780_));
 sky130_fd_sc_hd__o211a_1 _08754_ (.A1(_02778_),
    .A2(_02779_),
    .B1(_02613_),
    .C1(_02616_),
    .X(_02781_));
 sky130_fd_sc_hd__a22o_1 _08755_ (.A1(net200),
    .A2(net509),
    .B1(net502),
    .B2(net211),
    .X(_02782_));
 sky130_fd_sc_hd__and3_1 _08756_ (.A(net200),
    .B(net509),
    .C(net505),
    .X(_02783_));
 sky130_fd_sc_hd__and2_1 _08757_ (.A(net211),
    .B(_02783_),
    .X(_02784_));
 sky130_fd_sc_hd__a21bo_1 _08758_ (.A1(net211),
    .A2(_02783_),
    .B1_N(_02782_),
    .X(_02786_));
 sky130_fd_sc_hd__nand2_1 _08759_ (.A(net194),
    .B(net523),
    .Y(_02787_));
 sky130_fd_sc_hd__xor2_1 _08760_ (.A(_02786_),
    .B(_02787_),
    .X(_02788_));
 sky130_fd_sc_hd__and2_1 _08761_ (.A(_02649_),
    .B(_02653_),
    .X(_02789_));
 sky130_fd_sc_hd__and2b_1 _08762_ (.A_N(_02789_),
    .B(_02788_),
    .X(_02790_));
 sky130_fd_sc_hd__xor2_1 _08763_ (.A(_02788_),
    .B(_02789_),
    .X(_02791_));
 sky130_fd_sc_hd__or2_1 _08764_ (.A(_02659_),
    .B(_02791_),
    .X(_02792_));
 sky130_fd_sc_hd__xor2_1 _08765_ (.A(_02659_),
    .B(_02791_),
    .X(_02793_));
 sky130_fd_sc_hd__nand2_1 _08766_ (.A(_02637_),
    .B(_02639_),
    .Y(_02794_));
 sky130_fd_sc_hd__a21bo_1 _08767_ (.A1(_02646_),
    .A2(_02656_),
    .B1_N(_02655_),
    .X(_02795_));
 sky130_fd_sc_hd__and4_1 _08768_ (.A(net413),
    .B(net405),
    .C(net567),
    .D(net560),
    .X(_02797_));
 sky130_fd_sc_hd__a22o_1 _08769_ (.A1(net405),
    .A2(net567),
    .B1(net559),
    .B2(net413),
    .X(_02798_));
 sky130_fd_sc_hd__and2b_1 _08770_ (.A_N(_02797_),
    .B(_02798_),
    .X(_02799_));
 sky130_fd_sc_hd__nand2_1 _08771_ (.A(net398),
    .B(net574),
    .Y(_02800_));
 sky130_fd_sc_hd__xnor2_1 _08772_ (.A(_02799_),
    .B(_02800_),
    .Y(_02801_));
 sky130_fd_sc_hd__nand4_1 _08773_ (.A(net184),
    .B(net426),
    .C(net538),
    .D(net532),
    .Y(_02802_));
 sky130_fd_sc_hd__a22o_1 _08774_ (.A1(net426),
    .A2(net538),
    .B1(net532),
    .B2(net184),
    .X(_02803_));
 sky130_fd_sc_hd__and2_1 _08775_ (.A(net422),
    .B(net552),
    .X(_02804_));
 sky130_fd_sc_hd__a21o_1 _08776_ (.A1(_02802_),
    .A2(_02803_),
    .B1(_02804_),
    .X(_02805_));
 sky130_fd_sc_hd__nand3_1 _08777_ (.A(_02802_),
    .B(_02803_),
    .C(_02804_),
    .Y(_02806_));
 sky130_fd_sc_hd__a21bo_1 _08778_ (.A1(_02631_),
    .A2(_02633_),
    .B1_N(_02630_),
    .X(_02808_));
 sky130_fd_sc_hd__nand3_1 _08779_ (.A(_02805_),
    .B(_02806_),
    .C(_02808_),
    .Y(_02809_));
 sky130_fd_sc_hd__a21o_1 _08780_ (.A1(_02805_),
    .A2(_02806_),
    .B1(_02808_),
    .X(_02810_));
 sky130_fd_sc_hd__nand3_1 _08781_ (.A(_02801_),
    .B(_02809_),
    .C(_02810_),
    .Y(_02811_));
 sky130_fd_sc_hd__a21o_1 _08782_ (.A1(_02809_),
    .A2(_02810_),
    .B1(_02801_),
    .X(_02812_));
 sky130_fd_sc_hd__nand3_2 _08783_ (.A(_02795_),
    .B(_02811_),
    .C(_02812_),
    .Y(_02813_));
 sky130_fd_sc_hd__a21o_1 _08784_ (.A1(_02811_),
    .A2(_02812_),
    .B1(_02795_),
    .X(_02814_));
 sky130_fd_sc_hd__nand3_2 _08785_ (.A(_02794_),
    .B(_02813_),
    .C(_02814_),
    .Y(_02815_));
 sky130_fd_sc_hd__a21o_1 _08786_ (.A1(_02813_),
    .A2(_02814_),
    .B1(_02794_),
    .X(_02816_));
 sky130_fd_sc_hd__and3_1 _08787_ (.A(_02793_),
    .B(_02815_),
    .C(_02816_),
    .X(_02817_));
 sky130_fd_sc_hd__nand3_1 _08788_ (.A(_02793_),
    .B(_02815_),
    .C(_02816_),
    .Y(_02819_));
 sky130_fd_sc_hd__a21oi_1 _08789_ (.A1(_02815_),
    .A2(_02816_),
    .B1(_02793_),
    .Y(_02820_));
 sky130_fd_sc_hd__a211o_1 _08790_ (.A1(_02661_),
    .A2(_02663_),
    .B1(_02817_),
    .C1(_02820_),
    .X(_02821_));
 sky130_fd_sc_hd__o211ai_1 _08791_ (.A1(_02817_),
    .A2(_02820_),
    .B1(_02661_),
    .C1(_02663_),
    .Y(_02822_));
 sky130_fd_sc_hd__or4bb_2 _08792_ (.A(_02780_),
    .B(_02781_),
    .C_N(_02821_),
    .D_N(_02822_),
    .X(_02823_));
 sky130_fd_sc_hd__a2bb2o_1 _08793_ (.A1_N(_02780_),
    .A2_N(_02781_),
    .B1(_02821_),
    .B2(_02822_),
    .X(_02824_));
 sky130_fd_sc_hd__o211a_1 _08794_ (.A1(_02666_),
    .A2(net145),
    .B1(_02823_),
    .C1(_02824_),
    .X(_02825_));
 sky130_fd_sc_hd__a211oi_1 _08795_ (.A1(_02823_),
    .A2(_02824_),
    .B1(_02666_),
    .C1(net145),
    .Y(_02826_));
 sky130_fd_sc_hd__nor4_1 _08796_ (.A(_02740_),
    .B(_02742_),
    .C(_02825_),
    .D(_02826_),
    .Y(_02827_));
 sky130_fd_sc_hd__o22a_1 _08797_ (.A1(_02740_),
    .A2(_02742_),
    .B1(_02825_),
    .B2(_02826_),
    .X(_02828_));
 sky130_fd_sc_hd__nor2_1 _08798_ (.A(net135),
    .B(_02828_),
    .Y(_02830_));
 sky130_fd_sc_hd__a21boi_1 _08799_ (.A1(_02582_),
    .A2(_02673_),
    .B1_N(_02672_),
    .Y(_02831_));
 sky130_fd_sc_hd__and2b_1 _08800_ (.A_N(_02831_),
    .B(_02830_),
    .X(_02832_));
 sky130_fd_sc_hd__xnor2_1 _08801_ (.A(_02830_),
    .B(_02831_),
    .Y(_02833_));
 sky130_fd_sc_hd__xor2_1 _08802_ (.A(_02695_),
    .B(_02833_),
    .X(_02834_));
 sky130_fd_sc_hd__a21oi_1 _08803_ (.A1(_02537_),
    .A2(_02678_),
    .B1(_02677_),
    .Y(_02835_));
 sky130_fd_sc_hd__and2b_1 _08804_ (.A_N(_02835_),
    .B(_02834_),
    .X(_02836_));
 sky130_fd_sc_hd__xnor2_1 _08805_ (.A(_02834_),
    .B(_02835_),
    .Y(_02837_));
 sky130_fd_sc_hd__xnor2_1 _08806_ (.A(_02694_),
    .B(_02837_),
    .Y(_02838_));
 sky130_fd_sc_hd__a21o_1 _08807_ (.A1(_02682_),
    .A2(_02684_),
    .B1(_02838_),
    .X(_02839_));
 sky130_fd_sc_hd__inv_2 _08808_ (.A(_02839_),
    .Y(_02841_));
 sky130_fd_sc_hd__and3_1 _08809_ (.A(_02682_),
    .B(_02684_),
    .C(_02838_),
    .X(_02842_));
 sky130_fd_sc_hd__nor2_1 _08810_ (.A(_02841_),
    .B(_02842_),
    .Y(_02843_));
 sky130_fd_sc_hd__a21bo_1 _08811_ (.A1(_02689_),
    .A2(_02693_),
    .B1_N(_02688_),
    .X(_02844_));
 sky130_fd_sc_hd__xor2_1 _08812_ (.A(_02843_),
    .B(_02844_),
    .X(net95));
 sky130_fd_sc_hd__o21ai_1 _08813_ (.A1(_02706_),
    .A2(_02707_),
    .B1(_02711_),
    .Y(_02845_));
 sky130_fd_sc_hd__inv_2 _08814_ (.A(_02845_),
    .Y(_02846_));
 sky130_fd_sc_hd__nor2_1 _08815_ (.A(_02737_),
    .B(_02740_),
    .Y(_02847_));
 sky130_fd_sc_hd__and4_1 _08816_ (.A(net545),
    .B(net464),
    .C(net281),
    .D(net272),
    .X(_02848_));
 sky130_fd_sc_hd__a22oi_1 _08817_ (.A1(net464),
    .A2(net281),
    .B1(net272),
    .B2(net545),
    .Y(_02849_));
 sky130_fd_sc_hd__o2bb2a_1 _08818_ (.A1_N(net444),
    .A2_N(net263),
    .B1(_02848_),
    .B2(_02849_),
    .X(_02851_));
 sky130_fd_sc_hd__and4bb_1 _08819_ (.A_N(_02848_),
    .B_N(_02849_),
    .C(net444),
    .D(net263),
    .X(_02852_));
 sky130_fd_sc_hd__nor2_1 _08820_ (.A(_02851_),
    .B(_02852_),
    .Y(_02853_));
 sky130_fd_sc_hd__nor2_1 _08821_ (.A(_02696_),
    .B(_02700_),
    .Y(_02854_));
 sky130_fd_sc_hd__and2b_1 _08822_ (.A_N(_02854_),
    .B(_02853_),
    .X(_02855_));
 sky130_fd_sc_hd__xnor2_1 _08823_ (.A(_02853_),
    .B(_02854_),
    .Y(_02856_));
 sky130_fd_sc_hd__and2_1 _08824_ (.A(net31),
    .B(net252),
    .X(_02857_));
 sky130_fd_sc_hd__xnor2_1 _08825_ (.A(_02856_),
    .B(_02857_),
    .Y(_02858_));
 sky130_fd_sc_hd__a21oi_1 _08826_ (.A1(_02704_),
    .A2(_02705_),
    .B1(_02703_),
    .Y(_02859_));
 sky130_fd_sc_hd__xnor2_1 _08827_ (.A(_02858_),
    .B(_02859_),
    .Y(_02860_));
 sky130_fd_sc_hd__nand2_1 _08828_ (.A(net462),
    .B(net247),
    .Y(_02862_));
 sky130_fd_sc_hd__or2_1 _08829_ (.A(_02860_),
    .B(_02862_),
    .X(_02863_));
 sky130_fd_sc_hd__xor2_1 _08830_ (.A(_02860_),
    .B(_02862_),
    .X(_02864_));
 sky130_fd_sc_hd__a21o_1 _08831_ (.A1(_02747_),
    .A2(_02756_),
    .B1(_02755_),
    .X(_02865_));
 sky130_fd_sc_hd__nand2_1 _08832_ (.A(_02716_),
    .B(_02720_),
    .Y(_02866_));
 sky130_fd_sc_hd__a31o_1 _08833_ (.A1(net221),
    .A2(net313),
    .A3(_02744_),
    .B1(_02743_),
    .X(_02867_));
 sky130_fd_sc_hd__nand4_2 _08834_ (.A(net297),
    .B(net221),
    .C(net305),
    .D(net290),
    .Y(_02868_));
 sky130_fd_sc_hd__a22o_1 _08835_ (.A1(net221),
    .A2(net305),
    .B1(net290),
    .B2(net299),
    .X(_02869_));
 sky130_fd_sc_hd__a22o_1 _08836_ (.A1(net381),
    .A2(net283),
    .B1(_02868_),
    .B2(_02869_),
    .X(_02870_));
 sky130_fd_sc_hd__nand4_2 _08837_ (.A(net381),
    .B(net283),
    .C(_02868_),
    .D(_02869_),
    .Y(_02871_));
 sky130_fd_sc_hd__nand3_2 _08838_ (.A(_02867_),
    .B(_02870_),
    .C(_02871_),
    .Y(_02873_));
 sky130_fd_sc_hd__a21o_1 _08839_ (.A1(_02870_),
    .A2(_02871_),
    .B1(_02867_),
    .X(_02874_));
 sky130_fd_sc_hd__nand3_2 _08840_ (.A(_02866_),
    .B(_02873_),
    .C(_02874_),
    .Y(_02875_));
 sky130_fd_sc_hd__a21o_1 _08841_ (.A1(_02873_),
    .A2(_02874_),
    .B1(_02866_),
    .X(_02876_));
 sky130_fd_sc_hd__and3_2 _08842_ (.A(_02865_),
    .B(_02875_),
    .C(_02876_),
    .X(_02877_));
 sky130_fd_sc_hd__a21oi_2 _08843_ (.A1(_02875_),
    .A2(_02876_),
    .B1(_02865_),
    .Y(_02878_));
 sky130_fd_sc_hd__a211oi_2 _08844_ (.A1(_02721_),
    .A2(_02723_),
    .B1(_02877_),
    .C1(_02878_),
    .Y(_02879_));
 sky130_fd_sc_hd__a211o_1 _08845_ (.A1(_02721_),
    .A2(_02723_),
    .B1(_02877_),
    .C1(_02878_),
    .X(_02880_));
 sky130_fd_sc_hd__o211ai_2 _08846_ (.A1(_02877_),
    .A2(_02878_),
    .B1(_02721_),
    .C1(_02723_),
    .Y(_02881_));
 sky130_fd_sc_hd__o211ai_4 _08847_ (.A1(_02725_),
    .A2(_02727_),
    .B1(_02880_),
    .C1(_02881_),
    .Y(_02882_));
 sky130_fd_sc_hd__inv_2 _08848_ (.A(_02882_),
    .Y(_02884_));
 sky130_fd_sc_hd__a211o_1 _08849_ (.A1(_02880_),
    .A2(_02881_),
    .B1(_02725_),
    .C1(_02727_),
    .X(_02885_));
 sky130_fd_sc_hd__and3_1 _08850_ (.A(_02864_),
    .B(_02882_),
    .C(_02885_),
    .X(_02886_));
 sky130_fd_sc_hd__nand3_2 _08851_ (.A(_02864_),
    .B(_02882_),
    .C(_02885_),
    .Y(_02887_));
 sky130_fd_sc_hd__a21o_1 _08852_ (.A1(_02882_),
    .A2(_02885_),
    .B1(_02864_),
    .X(_02888_));
 sky130_fd_sc_hd__o211ai_4 _08853_ (.A1(_02778_),
    .A2(_02780_),
    .B1(_02887_),
    .C1(_02888_),
    .Y(_02889_));
 sky130_fd_sc_hd__a211o_1 _08854_ (.A1(_02887_),
    .A2(_02888_),
    .B1(_02778_),
    .C1(_02780_),
    .X(_02890_));
 sky130_fd_sc_hd__o211ai_4 _08855_ (.A1(_02732_),
    .A2(_02734_),
    .B1(_02889_),
    .C1(_02890_),
    .Y(_02891_));
 sky130_fd_sc_hd__a211o_1 _08856_ (.A1(_02889_),
    .A2(_02890_),
    .B1(_02732_),
    .C1(_02734_),
    .X(_02892_));
 sky130_fd_sc_hd__a22o_1 _08857_ (.A1(net194),
    .A2(net510),
    .B1(net503),
    .B2(net206),
    .X(_02893_));
 sky130_fd_sc_hd__nand2_1 _08858_ (.A(net194),
    .B(net503),
    .Y(_02895_));
 sky130_fd_sc_hd__o21a_1 _08859_ (.A1(_02648_),
    .A2(_02895_),
    .B1(_02893_),
    .X(_02896_));
 sky130_fd_sc_hd__a31o_1 _08860_ (.A1(net194),
    .A2(net524),
    .A3(_02782_),
    .B1(_02784_),
    .X(_02897_));
 sky130_fd_sc_hd__and2_1 _08861_ (.A(_02896_),
    .B(_02897_),
    .X(_02898_));
 sky130_fd_sc_hd__nor2_1 _08862_ (.A(_02896_),
    .B(_02897_),
    .Y(_02899_));
 sky130_fd_sc_hd__nor2_1 _08863_ (.A(_02898_),
    .B(_02899_),
    .Y(_02900_));
 sky130_fd_sc_hd__nand2_1 _08864_ (.A(_02809_),
    .B(_02811_),
    .Y(_02901_));
 sky130_fd_sc_hd__and4_1 _08865_ (.A(net413),
    .B(net405),
    .C(net560),
    .D(net553),
    .X(_02902_));
 sky130_fd_sc_hd__a22o_1 _08866_ (.A1(net405),
    .A2(net560),
    .B1(net553),
    .B2(net413),
    .X(_02903_));
 sky130_fd_sc_hd__and2b_1 _08867_ (.A_N(_02902_),
    .B(_02903_),
    .X(_02904_));
 sky130_fd_sc_hd__nand2_1 _08868_ (.A(net398),
    .B(net567),
    .Y(_02906_));
 sky130_fd_sc_hd__xnor2_1 _08869_ (.A(_02904_),
    .B(_02906_),
    .Y(_02907_));
 sky130_fd_sc_hd__nand4_1 _08870_ (.A(net186),
    .B(net426),
    .C(net532),
    .D(net523),
    .Y(_02908_));
 sky130_fd_sc_hd__a22o_1 _08871_ (.A1(net426),
    .A2(net532),
    .B1(net523),
    .B2(net186),
    .X(_02909_));
 sky130_fd_sc_hd__and2_1 _08872_ (.A(net422),
    .B(net539),
    .X(_02910_));
 sky130_fd_sc_hd__a21o_1 _08873_ (.A1(_02908_),
    .A2(_02909_),
    .B1(_02910_),
    .X(_02911_));
 sky130_fd_sc_hd__nand3_1 _08874_ (.A(_02908_),
    .B(_02909_),
    .C(_02910_),
    .Y(_02912_));
 sky130_fd_sc_hd__a21bo_1 _08875_ (.A1(_02803_),
    .A2(_02804_),
    .B1_N(_02802_),
    .X(_02913_));
 sky130_fd_sc_hd__nand3_1 _08876_ (.A(_02911_),
    .B(_02912_),
    .C(_02913_),
    .Y(_02914_));
 sky130_fd_sc_hd__a21o_1 _08877_ (.A1(_02911_),
    .A2(_02912_),
    .B1(_02913_),
    .X(_02915_));
 sky130_fd_sc_hd__nand3_1 _08878_ (.A(_02907_),
    .B(_02914_),
    .C(_02915_),
    .Y(_02917_));
 sky130_fd_sc_hd__a21o_1 _08879_ (.A1(_02914_),
    .A2(_02915_),
    .B1(_02907_),
    .X(_02918_));
 sky130_fd_sc_hd__nand3_2 _08880_ (.A(_02790_),
    .B(_02917_),
    .C(_02918_),
    .Y(_02919_));
 sky130_fd_sc_hd__a21o_1 _08881_ (.A1(_02917_),
    .A2(_02918_),
    .B1(_02790_),
    .X(_02920_));
 sky130_fd_sc_hd__nand3_2 _08882_ (.A(_02901_),
    .B(_02919_),
    .C(_02920_),
    .Y(_02921_));
 sky130_fd_sc_hd__a21o_1 _08883_ (.A1(_02919_),
    .A2(_02920_),
    .B1(_02901_),
    .X(_02922_));
 sky130_fd_sc_hd__and3_1 _08884_ (.A(_02900_),
    .B(_02921_),
    .C(_02922_),
    .X(_02923_));
 sky130_fd_sc_hd__a21oi_1 _08885_ (.A1(_02921_),
    .A2(_02922_),
    .B1(_02900_),
    .Y(_02924_));
 sky130_fd_sc_hd__o211a_1 _08886_ (.A1(_02923_),
    .A2(_02924_),
    .B1(_02792_),
    .C1(_02819_),
    .X(_02925_));
 sky130_fd_sc_hd__a211oi_2 _08887_ (.A1(_02792_),
    .A2(_02819_),
    .B1(_02923_),
    .C1(_02924_),
    .Y(_02926_));
 sky130_fd_sc_hd__inv_2 _08888_ (.A(_02926_),
    .Y(_02928_));
 sky130_fd_sc_hd__and4_1 _08889_ (.A(net169),
    .B(net161),
    .C(net328),
    .D(net320),
    .X(_02929_));
 sky130_fd_sc_hd__a22o_1 _08890_ (.A1(net161),
    .A2(net328),
    .B1(net320),
    .B2(net169),
    .X(_02930_));
 sky130_fd_sc_hd__and2b_1 _08891_ (.A_N(_02929_),
    .B(_02930_),
    .X(_02931_));
 sky130_fd_sc_hd__nand2_1 _08892_ (.A(net177),
    .B(net313),
    .Y(_02932_));
 sky130_fd_sc_hd__xnor2_1 _08893_ (.A(_02931_),
    .B(_02932_),
    .Y(_02933_));
 sky130_fd_sc_hd__nand4_1 _08894_ (.A(net358),
    .B(net611),
    .C(net350),
    .D(net595),
    .Y(_02934_));
 sky130_fd_sc_hd__a22o_1 _08895_ (.A1(net611),
    .A2(net350),
    .B1(net595),
    .B2(net358),
    .X(_02935_));
 sky130_fd_sc_hd__and2_1 _08896_ (.A(net623),
    .B(net335),
    .X(_02936_));
 sky130_fd_sc_hd__a21o_1 _08897_ (.A1(_02934_),
    .A2(_02935_),
    .B1(_02936_),
    .X(_02937_));
 sky130_fd_sc_hd__nand3_1 _08898_ (.A(_02934_),
    .B(_02935_),
    .C(_02936_),
    .Y(_02939_));
 sky130_fd_sc_hd__a21bo_1 _08899_ (.A1(_02749_),
    .A2(_02750_),
    .B1_N(_02748_),
    .X(_02940_));
 sky130_fd_sc_hd__and3_1 _08900_ (.A(_02937_),
    .B(_02939_),
    .C(_02940_),
    .X(_02941_));
 sky130_fd_sc_hd__a21o_1 _08901_ (.A1(_02937_),
    .A2(_02939_),
    .B1(_02940_),
    .X(_02942_));
 sky130_fd_sc_hd__and2b_1 _08902_ (.A_N(_02941_),
    .B(_02942_),
    .X(_02943_));
 sky130_fd_sc_hd__xnor2_1 _08903_ (.A(_02933_),
    .B(_02943_),
    .Y(_02944_));
 sky130_fd_sc_hd__nand2_1 _08904_ (.A(_02761_),
    .B(_02765_),
    .Y(_02945_));
 sky130_fd_sc_hd__a31o_1 _08905_ (.A1(net398),
    .A2(net574),
    .A3(_02798_),
    .B1(_02797_),
    .X(_02946_));
 sky130_fd_sc_hd__nand4_1 _08906_ (.A(net390),
    .B(net374),
    .C(net580),
    .D(net574),
    .Y(_02947_));
 sky130_fd_sc_hd__a22o_1 _08907_ (.A1(net374),
    .A2(net580),
    .B1(net574),
    .B2(net390),
    .X(_02948_));
 sky130_fd_sc_hd__a22o_1 _08908_ (.A1(net366),
    .A2(net588),
    .B1(_02947_),
    .B2(_02948_),
    .X(_02950_));
 sky130_fd_sc_hd__nand4_1 _08909_ (.A(net366),
    .B(net588),
    .C(_02947_),
    .D(_02948_),
    .Y(_02951_));
 sky130_fd_sc_hd__nand3_1 _08910_ (.A(_02946_),
    .B(_02950_),
    .C(_02951_),
    .Y(_02952_));
 sky130_fd_sc_hd__a21o_1 _08911_ (.A1(_02950_),
    .A2(_02951_),
    .B1(_02946_),
    .X(_02953_));
 sky130_fd_sc_hd__nand3_1 _08912_ (.A(_02945_),
    .B(_02952_),
    .C(_02953_),
    .Y(_02954_));
 sky130_fd_sc_hd__a21o_1 _08913_ (.A1(_02952_),
    .A2(_02953_),
    .B1(_02945_),
    .X(_02955_));
 sky130_fd_sc_hd__a21bo_1 _08914_ (.A1(_02759_),
    .A2(_02767_),
    .B1_N(_02766_),
    .X(_02956_));
 sky130_fd_sc_hd__and3_1 _08915_ (.A(_02954_),
    .B(_02955_),
    .C(_02956_),
    .X(_02957_));
 sky130_fd_sc_hd__inv_2 _08916_ (.A(_02957_),
    .Y(_02958_));
 sky130_fd_sc_hd__a21oi_1 _08917_ (.A1(_02954_),
    .A2(_02955_),
    .B1(_02956_),
    .Y(_02959_));
 sky130_fd_sc_hd__nor3_1 _08918_ (.A(_02944_),
    .B(_02957_),
    .C(_02959_),
    .Y(_02961_));
 sky130_fd_sc_hd__or3_1 _08919_ (.A(_02944_),
    .B(_02957_),
    .C(_02959_),
    .X(_02962_));
 sky130_fd_sc_hd__o21a_1 _08920_ (.A1(_02957_),
    .A2(_02959_),
    .B1(_02944_),
    .X(_02963_));
 sky130_fd_sc_hd__a211oi_4 _08921_ (.A1(_02813_),
    .A2(_02815_),
    .B1(net155),
    .C1(_02963_),
    .Y(_02964_));
 sky130_fd_sc_hd__o211a_1 _08922_ (.A1(_02961_),
    .A2(_02963_),
    .B1(_02813_),
    .C1(_02815_),
    .X(_02965_));
 sky130_fd_sc_hd__a211oi_4 _08923_ (.A1(_02772_),
    .A2(_02776_),
    .B1(_02964_),
    .C1(_02965_),
    .Y(_02966_));
 sky130_fd_sc_hd__o211a_1 _08924_ (.A1(_02964_),
    .A2(_02965_),
    .B1(_02772_),
    .C1(_02776_),
    .X(_02967_));
 sky130_fd_sc_hd__nor4_1 _08925_ (.A(_02925_),
    .B(_02926_),
    .C(_02966_),
    .D(_02967_),
    .Y(_02968_));
 sky130_fd_sc_hd__or4_1 _08926_ (.A(_02925_),
    .B(_02926_),
    .C(_02966_),
    .D(_02967_),
    .X(_02969_));
 sky130_fd_sc_hd__o22a_1 _08927_ (.A1(_02925_),
    .A2(_02926_),
    .B1(_02966_),
    .B2(_02967_),
    .X(_02970_));
 sky130_fd_sc_hd__a211o_2 _08928_ (.A1(_02821_),
    .A2(_02823_),
    .B1(_02968_),
    .C1(_02970_),
    .X(_02972_));
 sky130_fd_sc_hd__o211ai_2 _08929_ (.A1(net144),
    .A2(_02970_),
    .B1(_02821_),
    .C1(_02823_),
    .Y(_02973_));
 sky130_fd_sc_hd__nand4_4 _08930_ (.A(_02891_),
    .B(_02892_),
    .C(_02972_),
    .D(_02973_),
    .Y(_02974_));
 sky130_fd_sc_hd__a22o_1 _08931_ (.A1(_02891_),
    .A2(_02892_),
    .B1(_02972_),
    .B2(_02973_),
    .X(_02975_));
 sky130_fd_sc_hd__o211a_1 _08932_ (.A1(_02825_),
    .A2(_02827_),
    .B1(_02974_),
    .C1(_02975_),
    .X(_02976_));
 sky130_fd_sc_hd__a211oi_1 _08933_ (.A1(_02974_),
    .A2(_02975_),
    .B1(_02825_),
    .C1(net135),
    .Y(_02977_));
 sky130_fd_sc_hd__or3_1 _08934_ (.A(_02847_),
    .B(_02976_),
    .C(_02977_),
    .X(_02978_));
 sky130_fd_sc_hd__o21ai_1 _08935_ (.A1(_02976_),
    .A2(_02977_),
    .B1(_02847_),
    .Y(_02979_));
 sky130_fd_sc_hd__nand2_1 _08936_ (.A(_02978_),
    .B(_02979_),
    .Y(_02980_));
 sky130_fd_sc_hd__a21oi_1 _08937_ (.A1(_02695_),
    .A2(_02833_),
    .B1(_02832_),
    .Y(_02981_));
 sky130_fd_sc_hd__or2_1 _08938_ (.A(_02980_),
    .B(_02981_),
    .X(_02983_));
 sky130_fd_sc_hd__xnor2_1 _08939_ (.A(_02980_),
    .B(_02981_),
    .Y(_02984_));
 sky130_fd_sc_hd__xnor2_1 _08940_ (.A(_02846_),
    .B(_02984_),
    .Y(_02985_));
 sky130_fd_sc_hd__a21oi_1 _08941_ (.A1(_02694_),
    .A2(_02837_),
    .B1(_02836_),
    .Y(_02986_));
 sky130_fd_sc_hd__or2_1 _08942_ (.A(_02985_),
    .B(_02986_),
    .X(_02987_));
 sky130_fd_sc_hd__nand2_1 _08943_ (.A(_02985_),
    .B(_02986_),
    .Y(_02988_));
 sky130_fd_sc_hd__xnor2_1 _08944_ (.A(_02985_),
    .B(_02986_),
    .Y(_02989_));
 sky130_fd_sc_hd__a21oi_1 _08945_ (.A1(_02688_),
    .A2(_02839_),
    .B1(_02842_),
    .Y(_02990_));
 sky130_fd_sc_hd__and3b_1 _08946_ (.A_N(_02842_),
    .B(_02689_),
    .C(_02839_),
    .X(_02991_));
 sky130_fd_sc_hd__a21o_1 _08947_ (.A1(_02693_),
    .A2(_02991_),
    .B1(_02990_),
    .X(_02992_));
 sky130_fd_sc_hd__xnor2_1 _08948_ (.A(_02989_),
    .B(_02992_),
    .Y(net96));
 sky130_fd_sc_hd__o21a_1 _08949_ (.A1(_02858_),
    .A2(_02859_),
    .B1(_02863_),
    .X(_02994_));
 sky130_fd_sc_hd__nand2_1 _08950_ (.A(_02914_),
    .B(_02917_),
    .Y(_02995_));
 sky130_fd_sc_hd__and4_1 _08951_ (.A(net412),
    .B(net404),
    .C(net553),
    .D(net539),
    .X(_02996_));
 sky130_fd_sc_hd__a22o_1 _08952_ (.A1(net404),
    .A2(net553),
    .B1(net539),
    .B2(net412),
    .X(_02997_));
 sky130_fd_sc_hd__and2b_1 _08953_ (.A_N(_02996_),
    .B(_02997_),
    .X(_02998_));
 sky130_fd_sc_hd__nand2_1 _08954_ (.A(net398),
    .B(net560),
    .Y(_02999_));
 sky130_fd_sc_hd__xnor2_1 _08955_ (.A(_02998_),
    .B(_02999_),
    .Y(_03000_));
 sky130_fd_sc_hd__nand2_1 _08956_ (.A(net426),
    .B(net508),
    .Y(_03001_));
 sky130_fd_sc_hd__nand4_1 _08957_ (.A(net186),
    .B(net426),
    .C(net522),
    .D(net510),
    .Y(_03002_));
 sky130_fd_sc_hd__a22o_1 _08958_ (.A1(net433),
    .A2(net522),
    .B1(net510),
    .B2(net186),
    .X(_03004_));
 sky130_fd_sc_hd__and2_1 _08959_ (.A(net422),
    .B(net531),
    .X(_03005_));
 sky130_fd_sc_hd__a21o_1 _08960_ (.A1(_03002_),
    .A2(_03004_),
    .B1(_03005_),
    .X(_03006_));
 sky130_fd_sc_hd__nand3_1 _08961_ (.A(_03002_),
    .B(_03004_),
    .C(_03005_),
    .Y(_03007_));
 sky130_fd_sc_hd__a21bo_1 _08962_ (.A1(_02909_),
    .A2(_02910_),
    .B1_N(_02908_),
    .X(_03008_));
 sky130_fd_sc_hd__nand3_1 _08963_ (.A(_03006_),
    .B(_03007_),
    .C(_03008_),
    .Y(_03009_));
 sky130_fd_sc_hd__a21o_1 _08964_ (.A1(_03006_),
    .A2(_03007_),
    .B1(_03008_),
    .X(_03010_));
 sky130_fd_sc_hd__nand3_1 _08965_ (.A(_03000_),
    .B(_03009_),
    .C(_03010_),
    .Y(_03011_));
 sky130_fd_sc_hd__a21o_1 _08966_ (.A1(_03009_),
    .A2(_03010_),
    .B1(_03000_),
    .X(_03012_));
 sky130_fd_sc_hd__nand3_2 _08967_ (.A(_02898_),
    .B(_03011_),
    .C(_03012_),
    .Y(_03013_));
 sky130_fd_sc_hd__a21o_1 _08968_ (.A1(_03011_),
    .A2(_03012_),
    .B1(_02898_),
    .X(_03015_));
 sky130_fd_sc_hd__nand3_2 _08969_ (.A(_02995_),
    .B(_03013_),
    .C(_03015_),
    .Y(_03016_));
 sky130_fd_sc_hd__a21o_1 _08970_ (.A1(_03013_),
    .A2(_03015_),
    .B1(_02995_),
    .X(_03017_));
 sky130_fd_sc_hd__or4bb_2 _08971_ (.A(_02647_),
    .B(_02895_),
    .C_N(_03016_),
    .D_N(_03017_),
    .X(_03018_));
 sky130_fd_sc_hd__a2bb2o_1 _08972_ (.A1_N(_02647_),
    .A2_N(_02895_),
    .B1(_03016_),
    .B2(_03017_),
    .X(_03019_));
 sky130_fd_sc_hd__a21oi_1 _08973_ (.A1(_03018_),
    .A2(_03019_),
    .B1(_02923_),
    .Y(_03020_));
 sky130_fd_sc_hd__and3_1 _08974_ (.A(_02923_),
    .B(_03018_),
    .C(_03019_),
    .X(_03021_));
 sky130_fd_sc_hd__inv_2 _08975_ (.A(_03021_),
    .Y(_03022_));
 sky130_fd_sc_hd__and4_1 _08976_ (.A(net159),
    .B(net616),
    .C(net328),
    .D(net320),
    .X(_03023_));
 sky130_fd_sc_hd__a22o_1 _08977_ (.A1(net616),
    .A2(net328),
    .B1(net320),
    .B2(net159),
    .X(_03024_));
 sky130_fd_sc_hd__and2b_1 _08978_ (.A_N(_03023_),
    .B(_03024_),
    .X(_03026_));
 sky130_fd_sc_hd__nand2_1 _08979_ (.A(net168),
    .B(net313),
    .Y(_03027_));
 sky130_fd_sc_hd__xnor2_2 _08980_ (.A(_03026_),
    .B(_03027_),
    .Y(_03028_));
 sky130_fd_sc_hd__nand4_1 _08981_ (.A(net357),
    .B(net349),
    .C(net593),
    .D(net584),
    .Y(_03029_));
 sky130_fd_sc_hd__a22o_1 _08982_ (.A1(net349),
    .A2(net593),
    .B1(net586),
    .B2(net357),
    .X(_03030_));
 sky130_fd_sc_hd__and2_1 _08983_ (.A(net608),
    .B(net335),
    .X(_03031_));
 sky130_fd_sc_hd__a21o_1 _08984_ (.A1(_03029_),
    .A2(_03030_),
    .B1(_03031_),
    .X(_03032_));
 sky130_fd_sc_hd__nand3_1 _08985_ (.A(_03029_),
    .B(_03030_),
    .C(_03031_),
    .Y(_03033_));
 sky130_fd_sc_hd__a21bo_1 _08986_ (.A1(_02935_),
    .A2(_02936_),
    .B1_N(_02934_),
    .X(_03034_));
 sky130_fd_sc_hd__and3_1 _08987_ (.A(_03032_),
    .B(_03033_),
    .C(_03034_),
    .X(_03035_));
 sky130_fd_sc_hd__a21o_1 _08988_ (.A1(_03032_),
    .A2(_03033_),
    .B1(_03034_),
    .X(_03037_));
 sky130_fd_sc_hd__and2b_1 _08989_ (.A_N(_03035_),
    .B(_03037_),
    .X(_03038_));
 sky130_fd_sc_hd__xnor2_2 _08990_ (.A(_03028_),
    .B(_03038_),
    .Y(_03039_));
 sky130_fd_sc_hd__nand2_1 _08991_ (.A(_02947_),
    .B(_02951_),
    .Y(_03040_));
 sky130_fd_sc_hd__a31o_1 _08992_ (.A1(net398),
    .A2(net567),
    .A3(_02903_),
    .B1(_02902_),
    .X(_03041_));
 sky130_fd_sc_hd__nand4_1 _08993_ (.A(net389),
    .B(net373),
    .C(net574),
    .D(net567),
    .Y(_03042_));
 sky130_fd_sc_hd__a22o_1 _08994_ (.A1(net373),
    .A2(net574),
    .B1(net567),
    .B2(net389),
    .X(_03043_));
 sky130_fd_sc_hd__a22o_1 _08995_ (.A1(net366),
    .A2(net580),
    .B1(_03042_),
    .B2(_03043_),
    .X(_03044_));
 sky130_fd_sc_hd__nand4_1 _08996_ (.A(net366),
    .B(net580),
    .C(_03042_),
    .D(_03043_),
    .Y(_03045_));
 sky130_fd_sc_hd__nand3_1 _08997_ (.A(_03041_),
    .B(_03044_),
    .C(_03045_),
    .Y(_03046_));
 sky130_fd_sc_hd__a21o_1 _08998_ (.A1(_03044_),
    .A2(_03045_),
    .B1(_03041_),
    .X(_03048_));
 sky130_fd_sc_hd__nand3_1 _08999_ (.A(_03040_),
    .B(_03046_),
    .C(_03048_),
    .Y(_03049_));
 sky130_fd_sc_hd__a21o_1 _09000_ (.A1(_03046_),
    .A2(_03048_),
    .B1(_03040_),
    .X(_03050_));
 sky130_fd_sc_hd__a21bo_1 _09001_ (.A1(_02945_),
    .A2(_02953_),
    .B1_N(_02952_),
    .X(_03051_));
 sky130_fd_sc_hd__and3_2 _09002_ (.A(_03049_),
    .B(_03050_),
    .C(_03051_),
    .X(_03052_));
 sky130_fd_sc_hd__a21oi_2 _09003_ (.A1(_03049_),
    .A2(_03050_),
    .B1(_03051_),
    .Y(_03053_));
 sky130_fd_sc_hd__nor3_4 _09004_ (.A(_03039_),
    .B(_03052_),
    .C(_03053_),
    .Y(_03054_));
 sky130_fd_sc_hd__o21a_1 _09005_ (.A1(_03052_),
    .A2(_03053_),
    .B1(_03039_),
    .X(_03055_));
 sky130_fd_sc_hd__a211oi_4 _09006_ (.A1(_02919_),
    .A2(_02921_),
    .B1(_03054_),
    .C1(_03055_),
    .Y(_03056_));
 sky130_fd_sc_hd__o211a_1 _09007_ (.A1(_03054_),
    .A2(_03055_),
    .B1(_02919_),
    .C1(_02921_),
    .X(_03057_));
 sky130_fd_sc_hd__a211oi_2 _09008_ (.A1(_02958_),
    .A2(_02962_),
    .B1(_03056_),
    .C1(_03057_),
    .Y(_03059_));
 sky130_fd_sc_hd__o211a_1 _09009_ (.A1(_03056_),
    .A2(_03057_),
    .B1(_02958_),
    .C1(_02962_),
    .X(_03060_));
 sky130_fd_sc_hd__nor4_1 _09010_ (.A(_03020_),
    .B(_03021_),
    .C(_03059_),
    .D(_03060_),
    .Y(_03061_));
 sky130_fd_sc_hd__or4_1 _09011_ (.A(_03020_),
    .B(_03021_),
    .C(_03059_),
    .D(_03060_),
    .X(_03062_));
 sky130_fd_sc_hd__o22a_1 _09012_ (.A1(_03020_),
    .A2(_03021_),
    .B1(_03059_),
    .B2(_03060_),
    .X(_03063_));
 sky130_fd_sc_hd__a211oi_2 _09013_ (.A1(_02928_),
    .A2(_02969_),
    .B1(net143),
    .C1(_03063_),
    .Y(_03064_));
 sky130_fd_sc_hd__inv_2 _09014_ (.A(_03064_),
    .Y(_03065_));
 sky130_fd_sc_hd__o211a_1 _09015_ (.A1(_03061_),
    .A2(_03063_),
    .B1(_02928_),
    .C1(_02969_),
    .X(_03066_));
 sky130_fd_sc_hd__and4_1 _09016_ (.A(net464),
    .B(net381),
    .C(net276),
    .D(net268),
    .X(_03067_));
 sky130_fd_sc_hd__a22oi_1 _09017_ (.A1(net383),
    .A2(net276),
    .B1(net268),
    .B2(net464),
    .Y(_03068_));
 sky130_fd_sc_hd__o2bb2a_1 _09018_ (.A1_N(net545),
    .A2_N(net260),
    .B1(_03067_),
    .B2(_03068_),
    .X(_03070_));
 sky130_fd_sc_hd__and4bb_1 _09019_ (.A_N(_03067_),
    .B_N(_03068_),
    .C(net545),
    .D(net260),
    .X(_03071_));
 sky130_fd_sc_hd__nor2_1 _09020_ (.A(_03070_),
    .B(_03071_),
    .Y(_03072_));
 sky130_fd_sc_hd__nor2_1 _09021_ (.A(_02848_),
    .B(_02852_),
    .Y(_03073_));
 sky130_fd_sc_hd__or3_1 _09022_ (.A(_03070_),
    .B(_03071_),
    .C(_03073_),
    .X(_03074_));
 sky130_fd_sc_hd__xnor2_1 _09023_ (.A(_03072_),
    .B(_03073_),
    .Y(_03075_));
 sky130_fd_sc_hd__nand2_1 _09024_ (.A(net444),
    .B(net252),
    .Y(_03076_));
 sky130_fd_sc_hd__nand3_1 _09025_ (.A(net444),
    .B(net252),
    .C(_03075_),
    .Y(_03077_));
 sky130_fd_sc_hd__xor2_1 _09026_ (.A(_03075_),
    .B(_03076_),
    .X(_03078_));
 sky130_fd_sc_hd__a21oi_1 _09027_ (.A1(_02856_),
    .A2(_02857_),
    .B1(_02855_),
    .Y(_03079_));
 sky130_fd_sc_hd__xnor2_1 _09028_ (.A(_03078_),
    .B(_03079_),
    .Y(_03081_));
 sky130_fd_sc_hd__nand2_1 _09029_ (.A(net31),
    .B(net247),
    .Y(_03082_));
 sky130_fd_sc_hd__or2_1 _09030_ (.A(_03081_),
    .B(_03082_),
    .X(_03083_));
 sky130_fd_sc_hd__xor2_1 _09031_ (.A(_03081_),
    .B(_03082_),
    .X(_03084_));
 sky130_fd_sc_hd__a21o_1 _09032_ (.A1(_02933_),
    .A2(_02942_),
    .B1(_02941_),
    .X(_03085_));
 sky130_fd_sc_hd__nand2_1 _09033_ (.A(_02868_),
    .B(_02871_),
    .Y(_03086_));
 sky130_fd_sc_hd__a31o_1 _09034_ (.A1(net177),
    .A2(net313),
    .A3(_02930_),
    .B1(_02929_),
    .X(_03087_));
 sky130_fd_sc_hd__nand4_2 _09035_ (.A(net220),
    .B(net175),
    .C(net305),
    .D(net293),
    .Y(_03088_));
 sky130_fd_sc_hd__a22o_1 _09036_ (.A1(net176),
    .A2(net305),
    .B1(net293),
    .B2(net220),
    .X(_03089_));
 sky130_fd_sc_hd__a22o_1 _09037_ (.A1(net299),
    .A2(net286),
    .B1(_03088_),
    .B2(_03089_),
    .X(_03090_));
 sky130_fd_sc_hd__nand4_2 _09038_ (.A(net299),
    .B(net286),
    .C(_03088_),
    .D(_03089_),
    .Y(_03092_));
 sky130_fd_sc_hd__nand3_2 _09039_ (.A(_03087_),
    .B(_03090_),
    .C(_03092_),
    .Y(_03093_));
 sky130_fd_sc_hd__a21o_1 _09040_ (.A1(_03090_),
    .A2(_03092_),
    .B1(_03087_),
    .X(_03094_));
 sky130_fd_sc_hd__nand3_2 _09041_ (.A(_03086_),
    .B(_03093_),
    .C(_03094_),
    .Y(_03095_));
 sky130_fd_sc_hd__a21o_1 _09042_ (.A1(_03093_),
    .A2(_03094_),
    .B1(_03086_),
    .X(_03096_));
 sky130_fd_sc_hd__and3_2 _09043_ (.A(_03085_),
    .B(_03095_),
    .C(_03096_),
    .X(_03097_));
 sky130_fd_sc_hd__a21oi_2 _09044_ (.A1(_03095_),
    .A2(_03096_),
    .B1(_03085_),
    .Y(_03098_));
 sky130_fd_sc_hd__a211oi_2 _09045_ (.A1(_02873_),
    .A2(_02875_),
    .B1(_03097_),
    .C1(_03098_),
    .Y(_03099_));
 sky130_fd_sc_hd__a211o_1 _09046_ (.A1(_02873_),
    .A2(_02875_),
    .B1(_03097_),
    .C1(_03098_),
    .X(_03100_));
 sky130_fd_sc_hd__o211ai_2 _09047_ (.A1(_03097_),
    .A2(_03098_),
    .B1(_02873_),
    .C1(_02875_),
    .Y(_03101_));
 sky130_fd_sc_hd__o211ai_2 _09048_ (.A1(_02877_),
    .A2(_02879_),
    .B1(_03100_),
    .C1(_03101_),
    .Y(_03103_));
 sky130_fd_sc_hd__a211o_1 _09049_ (.A1(_03100_),
    .A2(_03101_),
    .B1(_02877_),
    .C1(_02879_),
    .X(_03104_));
 sky130_fd_sc_hd__nand3_2 _09050_ (.A(_03084_),
    .B(_03103_),
    .C(_03104_),
    .Y(_03105_));
 sky130_fd_sc_hd__a21o_1 _09051_ (.A1(_03103_),
    .A2(_03104_),
    .B1(_03084_),
    .X(_03106_));
 sky130_fd_sc_hd__o211ai_4 _09052_ (.A1(_02964_),
    .A2(_02966_),
    .B1(_03105_),
    .C1(_03106_),
    .Y(_03107_));
 sky130_fd_sc_hd__a211o_1 _09053_ (.A1(_03105_),
    .A2(_03106_),
    .B1(_02964_),
    .C1(_02966_),
    .X(_03108_));
 sky130_fd_sc_hd__o211ai_4 _09054_ (.A1(_02884_),
    .A2(_02886_),
    .B1(_03107_),
    .C1(_03108_),
    .Y(_03109_));
 sky130_fd_sc_hd__a211o_1 _09055_ (.A1(_03107_),
    .A2(_03108_),
    .B1(_02884_),
    .C1(_02886_),
    .X(_03110_));
 sky130_fd_sc_hd__and4bb_1 _09056_ (.A_N(_03064_),
    .B_N(_03066_),
    .C(_03109_),
    .D(_03110_),
    .X(_03111_));
 sky130_fd_sc_hd__or4bb_1 _09057_ (.A(_03064_),
    .B(_03066_),
    .C_N(_03109_),
    .D_N(_03110_),
    .X(_03112_));
 sky130_fd_sc_hd__a2bb2oi_2 _09058_ (.A1_N(_03064_),
    .A2_N(_03066_),
    .B1(_03109_),
    .B2(_03110_),
    .Y(_03114_));
 sky130_fd_sc_hd__a211oi_4 _09059_ (.A1(_02972_),
    .A2(_02974_),
    .B1(_03111_),
    .C1(_03114_),
    .Y(_03115_));
 sky130_fd_sc_hd__o211a_1 _09060_ (.A1(_03111_),
    .A2(_03114_),
    .B1(_02972_),
    .C1(_02974_),
    .X(_03116_));
 sky130_fd_sc_hd__a211oi_2 _09061_ (.A1(_02889_),
    .A2(_02891_),
    .B1(_03115_),
    .C1(_03116_),
    .Y(_03117_));
 sky130_fd_sc_hd__o211a_1 _09062_ (.A1(_03115_),
    .A2(_03116_),
    .B1(_02889_),
    .C1(_02891_),
    .X(_03118_));
 sky130_fd_sc_hd__o21ba_1 _09063_ (.A1(_02847_),
    .A2(_02977_),
    .B1_N(_02976_),
    .X(_03119_));
 sky130_fd_sc_hd__nor3_1 _09064_ (.A(_03117_),
    .B(_03118_),
    .C(_03119_),
    .Y(_03120_));
 sky130_fd_sc_hd__o21a_1 _09065_ (.A1(_03117_),
    .A2(_03118_),
    .B1(_03119_),
    .X(_03121_));
 sky130_fd_sc_hd__nor3_1 _09066_ (.A(_02994_),
    .B(net129),
    .C(_03121_),
    .Y(_03122_));
 sky130_fd_sc_hd__o21a_1 _09067_ (.A1(_03120_),
    .A2(_03121_),
    .B1(_02994_),
    .X(_03123_));
 sky130_fd_sc_hd__or2_1 _09068_ (.A(_03122_),
    .B(_03123_),
    .X(_03125_));
 sky130_fd_sc_hd__o21a_1 _09069_ (.A1(_02846_),
    .A2(_02984_),
    .B1(_02983_),
    .X(_03126_));
 sky130_fd_sc_hd__xnor2_1 _09070_ (.A(_03125_),
    .B(_03126_),
    .Y(_03127_));
 sky130_fd_sc_hd__a21bo_1 _09071_ (.A1(_02988_),
    .A2(_02992_),
    .B1_N(_02987_),
    .X(_03128_));
 sky130_fd_sc_hd__xnor2_1 _09072_ (.A(_03127_),
    .B(_03128_),
    .Y(net97));
 sky130_fd_sc_hd__o21ai_1 _09073_ (.A1(_03078_),
    .A2(_03079_),
    .B1(_03083_),
    .Y(_03129_));
 sky130_fd_sc_hd__and4_1 _09074_ (.A(net412),
    .B(net404),
    .C(net539),
    .D(net531),
    .X(_03130_));
 sky130_fd_sc_hd__a22o_1 _09075_ (.A1(net405),
    .A2(net539),
    .B1(net531),
    .B2(net412),
    .X(_03131_));
 sky130_fd_sc_hd__and2b_1 _09076_ (.A_N(_03130_),
    .B(_03131_),
    .X(_03132_));
 sky130_fd_sc_hd__nand2_1 _09077_ (.A(net397),
    .B(net553),
    .Y(_03133_));
 sky130_fd_sc_hd__xnor2_1 _09078_ (.A(_03132_),
    .B(_03133_),
    .Y(_03135_));
 sky130_fd_sc_hd__nand4_2 _09079_ (.A(net186),
    .B(net426),
    .C(net508),
    .D(net503),
    .Y(_03136_));
 sky130_fd_sc_hd__a22o_1 _09080_ (.A1(net426),
    .A2(net508),
    .B1(net503),
    .B2(net186),
    .X(_03137_));
 sky130_fd_sc_hd__a22o_1 _09081_ (.A1(net422),
    .A2(net522),
    .B1(_03136_),
    .B2(_03137_),
    .X(_03138_));
 sky130_fd_sc_hd__nand4_2 _09082_ (.A(net422),
    .B(net522),
    .C(_03136_),
    .D(_03137_),
    .Y(_03139_));
 sky130_fd_sc_hd__a21bo_1 _09083_ (.A1(_03004_),
    .A2(_03005_),
    .B1_N(_03002_),
    .X(_03140_));
 sky130_fd_sc_hd__and3_1 _09084_ (.A(_03138_),
    .B(_03139_),
    .C(_03140_),
    .X(_03141_));
 sky130_fd_sc_hd__a21oi_1 _09085_ (.A1(_03138_),
    .A2(_03139_),
    .B1(_03140_),
    .Y(_03142_));
 sky130_fd_sc_hd__nor3b_1 _09086_ (.A(_03141_),
    .B(_03142_),
    .C_N(_03135_),
    .Y(_03143_));
 sky130_fd_sc_hd__or3b_1 _09087_ (.A(_03141_),
    .B(_03142_),
    .C_N(_03135_),
    .X(_03144_));
 sky130_fd_sc_hd__o21bai_1 _09088_ (.A1(_03141_),
    .A2(_03142_),
    .B1_N(_03135_),
    .Y(_03146_));
 sky130_fd_sc_hd__or4b_2 _09089_ (.A(_02648_),
    .B(_02895_),
    .C(_03143_),
    .D_N(_03146_),
    .X(_03147_));
 sky130_fd_sc_hd__a2bb2o_1 _09090_ (.A1_N(_02648_),
    .A2_N(_02895_),
    .B1(_03144_),
    .B2(_03146_),
    .X(_03148_));
 sky130_fd_sc_hd__nand2_1 _09091_ (.A(_03009_),
    .B(_03011_),
    .Y(_03149_));
 sky130_fd_sc_hd__a21o_1 _09092_ (.A1(_03147_),
    .A2(_03148_),
    .B1(_03149_),
    .X(_03150_));
 sky130_fd_sc_hd__nand3_1 _09093_ (.A(_03147_),
    .B(_03148_),
    .C(_03149_),
    .Y(_03151_));
 sky130_fd_sc_hd__nand2_1 _09094_ (.A(_03150_),
    .B(_03151_),
    .Y(_03152_));
 sky130_fd_sc_hd__nor2_1 _09095_ (.A(_03018_),
    .B(_03152_),
    .Y(_03153_));
 sky130_fd_sc_hd__xor2_1 _09096_ (.A(_03018_),
    .B(_03152_),
    .X(_03154_));
 sky130_fd_sc_hd__and4_1 _09097_ (.A(net616),
    .B(net608),
    .C(net327),
    .D(net319),
    .X(_03155_));
 sky130_fd_sc_hd__a22o_1 _09098_ (.A1(net608),
    .A2(net327),
    .B1(net319),
    .B2(net616),
    .X(_03157_));
 sky130_fd_sc_hd__and2b_1 _09099_ (.A_N(_03155_),
    .B(_03157_),
    .X(_03158_));
 sky130_fd_sc_hd__nand2_1 _09100_ (.A(net160),
    .B(net312),
    .Y(_03159_));
 sky130_fd_sc_hd__xnor2_1 _09101_ (.A(_03158_),
    .B(_03159_),
    .Y(_03160_));
 sky130_fd_sc_hd__nand4_1 _09102_ (.A(net357),
    .B(net349),
    .C(net586),
    .D(net577),
    .Y(_03161_));
 sky130_fd_sc_hd__a22o_1 _09103_ (.A1(net349),
    .A2(net586),
    .B1(net578),
    .B2(net357),
    .X(_03162_));
 sky130_fd_sc_hd__and2_1 _09104_ (.A(net593),
    .B(net335),
    .X(_03163_));
 sky130_fd_sc_hd__a21o_1 _09105_ (.A1(_03161_),
    .A2(_03162_),
    .B1(_03163_),
    .X(_03164_));
 sky130_fd_sc_hd__nand3_1 _09106_ (.A(_03161_),
    .B(_03162_),
    .C(_03163_),
    .Y(_03165_));
 sky130_fd_sc_hd__a21bo_1 _09107_ (.A1(_03030_),
    .A2(_03031_),
    .B1_N(_03029_),
    .X(_03166_));
 sky130_fd_sc_hd__and3_1 _09108_ (.A(_03164_),
    .B(_03165_),
    .C(_03166_),
    .X(_03168_));
 sky130_fd_sc_hd__a21o_1 _09109_ (.A1(_03164_),
    .A2(_03165_),
    .B1(_03166_),
    .X(_03169_));
 sky130_fd_sc_hd__and2b_1 _09110_ (.A_N(_03168_),
    .B(_03169_),
    .X(_03170_));
 sky130_fd_sc_hd__xnor2_1 _09111_ (.A(_03160_),
    .B(_03170_),
    .Y(_03171_));
 sky130_fd_sc_hd__nand2_1 _09112_ (.A(_03042_),
    .B(_03045_),
    .Y(_03172_));
 sky130_fd_sc_hd__a31o_1 _09113_ (.A1(net398),
    .A2(net560),
    .A3(_02997_),
    .B1(_02996_),
    .X(_03173_));
 sky130_fd_sc_hd__nand4_1 _09114_ (.A(net389),
    .B(net373),
    .C(net567),
    .D(net560),
    .Y(_03174_));
 sky130_fd_sc_hd__a22o_1 _09115_ (.A1(net373),
    .A2(net567),
    .B1(net560),
    .B2(net389),
    .X(_03175_));
 sky130_fd_sc_hd__a22o_1 _09116_ (.A1(net365),
    .A2(net571),
    .B1(_03174_),
    .B2(_03175_),
    .X(_03176_));
 sky130_fd_sc_hd__nand4_1 _09117_ (.A(net365),
    .B(net572),
    .C(_03174_),
    .D(_03175_),
    .Y(_03177_));
 sky130_fd_sc_hd__nand3_1 _09118_ (.A(_03173_),
    .B(_03176_),
    .C(_03177_),
    .Y(_03179_));
 sky130_fd_sc_hd__a21o_1 _09119_ (.A1(_03176_),
    .A2(_03177_),
    .B1(_03173_),
    .X(_03180_));
 sky130_fd_sc_hd__nand3_1 _09120_ (.A(_03172_),
    .B(_03179_),
    .C(_03180_),
    .Y(_03181_));
 sky130_fd_sc_hd__a21o_1 _09121_ (.A1(_03179_),
    .A2(_03180_),
    .B1(_03172_),
    .X(_03182_));
 sky130_fd_sc_hd__a21bo_1 _09122_ (.A1(_03040_),
    .A2(_03048_),
    .B1_N(_03046_),
    .X(_03183_));
 sky130_fd_sc_hd__and3_1 _09123_ (.A(_03181_),
    .B(_03182_),
    .C(_03183_),
    .X(_03184_));
 sky130_fd_sc_hd__inv_2 _09124_ (.A(_03184_),
    .Y(_03185_));
 sky130_fd_sc_hd__a21oi_1 _09125_ (.A1(_03181_),
    .A2(_03182_),
    .B1(_03183_),
    .Y(_03186_));
 sky130_fd_sc_hd__nor3_1 _09126_ (.A(_03171_),
    .B(_03184_),
    .C(_03186_),
    .Y(_03187_));
 sky130_fd_sc_hd__inv_2 _09127_ (.A(_03187_),
    .Y(_03188_));
 sky130_fd_sc_hd__o21a_1 _09128_ (.A1(_03184_),
    .A2(_03186_),
    .B1(_03171_),
    .X(_03190_));
 sky130_fd_sc_hd__a211o_2 _09129_ (.A1(_03013_),
    .A2(_03016_),
    .B1(net154),
    .C1(_03190_),
    .X(_03191_));
 sky130_fd_sc_hd__o211ai_2 _09130_ (.A1(net154),
    .A2(_03190_),
    .B1(_03013_),
    .C1(_03016_),
    .Y(_03192_));
 sky130_fd_sc_hd__o211ai_4 _09131_ (.A1(_03052_),
    .A2(_03054_),
    .B1(_03191_),
    .C1(_03192_),
    .Y(_03193_));
 sky130_fd_sc_hd__a211o_1 _09132_ (.A1(_03191_),
    .A2(_03192_),
    .B1(_03052_),
    .C1(_03054_),
    .X(_03194_));
 sky130_fd_sc_hd__and3_2 _09133_ (.A(_03154_),
    .B(_03193_),
    .C(_03194_),
    .X(_03195_));
 sky130_fd_sc_hd__a21oi_1 _09134_ (.A1(_03193_),
    .A2(_03194_),
    .B1(_03154_),
    .Y(_03196_));
 sky130_fd_sc_hd__a211oi_2 _09135_ (.A1(_03022_),
    .A2(_03062_),
    .B1(_03195_),
    .C1(_03196_),
    .Y(_03197_));
 sky130_fd_sc_hd__o211a_1 _09136_ (.A1(_03195_),
    .A2(_03196_),
    .B1(_03022_),
    .C1(_03062_),
    .X(_03198_));
 sky130_fd_sc_hd__nand2_1 _09137_ (.A(_03103_),
    .B(_03105_),
    .Y(_03199_));
 sky130_fd_sc_hd__and4_1 _09138_ (.A(net381),
    .B(net297),
    .C(net276),
    .D(net268),
    .X(_03201_));
 sky130_fd_sc_hd__a22oi_1 _09139_ (.A1(net297),
    .A2(net276),
    .B1(net268),
    .B2(net381),
    .Y(_03202_));
 sky130_fd_sc_hd__o2bb2a_1 _09140_ (.A1_N(net464),
    .A2_N(net260),
    .B1(_03201_),
    .B2(_03202_),
    .X(_03203_));
 sky130_fd_sc_hd__and4bb_1 _09141_ (.A_N(_03201_),
    .B_N(_03202_),
    .C(net464),
    .D(net260),
    .X(_03204_));
 sky130_fd_sc_hd__nor2_1 _09142_ (.A(_03203_),
    .B(_03204_),
    .Y(_03205_));
 sky130_fd_sc_hd__nor2_1 _09143_ (.A(_03067_),
    .B(_03071_),
    .Y(_03206_));
 sky130_fd_sc_hd__and2b_1 _09144_ (.A_N(_03206_),
    .B(_03205_),
    .X(_03207_));
 sky130_fd_sc_hd__xnor2_1 _09145_ (.A(_03205_),
    .B(_03206_),
    .Y(_03208_));
 sky130_fd_sc_hd__and2_1 _09146_ (.A(net545),
    .B(net249),
    .X(_03209_));
 sky130_fd_sc_hd__xnor2_1 _09147_ (.A(_03208_),
    .B(_03209_),
    .Y(_03210_));
 sky130_fd_sc_hd__and3_1 _09148_ (.A(_03074_),
    .B(_03077_),
    .C(_03210_),
    .X(_03212_));
 sky130_fd_sc_hd__a21o_1 _09149_ (.A1(_03074_),
    .A2(_03077_),
    .B1(_03210_),
    .X(_03213_));
 sky130_fd_sc_hd__and2b_1 _09150_ (.A_N(_03212_),
    .B(_03213_),
    .X(_03214_));
 sky130_fd_sc_hd__nand2_1 _09151_ (.A(net444),
    .B(net243),
    .Y(_03215_));
 sky130_fd_sc_hd__nand3_1 _09152_ (.A(net444),
    .B(net246),
    .C(_03214_),
    .Y(_03216_));
 sky130_fd_sc_hd__xnor2_1 _09153_ (.A(_03214_),
    .B(_03215_),
    .Y(_03217_));
 sky130_fd_sc_hd__a21o_1 _09154_ (.A1(_03028_),
    .A2(_03037_),
    .B1(_03035_),
    .X(_03218_));
 sky130_fd_sc_hd__nand2_1 _09155_ (.A(_03088_),
    .B(_03092_),
    .Y(_03219_));
 sky130_fd_sc_hd__a31o_1 _09156_ (.A1(net168),
    .A2(net313),
    .A3(_03024_),
    .B1(_03023_),
    .X(_03220_));
 sky130_fd_sc_hd__nand4_2 _09157_ (.A(net176),
    .B(net168),
    .C(net304),
    .D(net293),
    .Y(_03221_));
 sky130_fd_sc_hd__a22o_1 _09158_ (.A1(net168),
    .A2(net305),
    .B1(net293),
    .B2(net176),
    .X(_03223_));
 sky130_fd_sc_hd__a22o_1 _09159_ (.A1(net223),
    .A2(net286),
    .B1(_03221_),
    .B2(_03223_),
    .X(_03224_));
 sky130_fd_sc_hd__nand4_2 _09160_ (.A(net223),
    .B(net286),
    .C(_03221_),
    .D(_03223_),
    .Y(_03225_));
 sky130_fd_sc_hd__nand3_2 _09161_ (.A(_03220_),
    .B(_03224_),
    .C(_03225_),
    .Y(_03226_));
 sky130_fd_sc_hd__a21o_1 _09162_ (.A1(_03224_),
    .A2(_03225_),
    .B1(_03220_),
    .X(_03227_));
 sky130_fd_sc_hd__nand3_2 _09163_ (.A(_03219_),
    .B(_03226_),
    .C(_03227_),
    .Y(_03228_));
 sky130_fd_sc_hd__a21o_1 _09164_ (.A1(_03226_),
    .A2(_03227_),
    .B1(_03219_),
    .X(_03229_));
 sky130_fd_sc_hd__and3_1 _09165_ (.A(_03218_),
    .B(_03228_),
    .C(_03229_),
    .X(_03230_));
 sky130_fd_sc_hd__nand3_1 _09166_ (.A(_03218_),
    .B(_03228_),
    .C(_03229_),
    .Y(_03231_));
 sky130_fd_sc_hd__a21oi_1 _09167_ (.A1(_03228_),
    .A2(_03229_),
    .B1(_03218_),
    .Y(_03232_));
 sky130_fd_sc_hd__a211o_2 _09168_ (.A1(_03093_),
    .A2(_03095_),
    .B1(_03230_),
    .C1(_03232_),
    .X(_03234_));
 sky130_fd_sc_hd__o211ai_2 _09169_ (.A1(_03230_),
    .A2(_03232_),
    .B1(_03093_),
    .C1(_03095_),
    .Y(_03235_));
 sky130_fd_sc_hd__o211ai_4 _09170_ (.A1(_03097_),
    .A2(_03099_),
    .B1(_03234_),
    .C1(_03235_),
    .Y(_03236_));
 sky130_fd_sc_hd__a211o_1 _09171_ (.A1(_03234_),
    .A2(_03235_),
    .B1(_03097_),
    .C1(_03099_),
    .X(_03237_));
 sky130_fd_sc_hd__nand3_2 _09172_ (.A(_03217_),
    .B(_03236_),
    .C(_03237_),
    .Y(_03238_));
 sky130_fd_sc_hd__a21o_1 _09173_ (.A1(_03236_),
    .A2(_03237_),
    .B1(_03217_),
    .X(_03239_));
 sky130_fd_sc_hd__o211ai_2 _09174_ (.A1(_03056_),
    .A2(_03059_),
    .B1(_03238_),
    .C1(_03239_),
    .Y(_03240_));
 sky130_fd_sc_hd__a211o_1 _09175_ (.A1(_03238_),
    .A2(_03239_),
    .B1(_03056_),
    .C1(_03059_),
    .X(_03241_));
 sky130_fd_sc_hd__nand3_1 _09176_ (.A(_03199_),
    .B(_03240_),
    .C(_03241_),
    .Y(_03242_));
 sky130_fd_sc_hd__a21o_1 _09177_ (.A1(_03240_),
    .A2(_03241_),
    .B1(_03199_),
    .X(_03243_));
 sky130_fd_sc_hd__and4bb_1 _09178_ (.A_N(_03197_),
    .B_N(_03198_),
    .C(_03242_),
    .D(_03243_),
    .X(_03245_));
 sky130_fd_sc_hd__a2bb2oi_1 _09179_ (.A1_N(_03197_),
    .A2_N(_03198_),
    .B1(_03242_),
    .B2(_03243_),
    .Y(_03246_));
 sky130_fd_sc_hd__a211oi_1 _09180_ (.A1(_03065_),
    .A2(_03112_),
    .B1(_03245_),
    .C1(_03246_),
    .Y(_03247_));
 sky130_fd_sc_hd__a211o_1 _09181_ (.A1(_03065_),
    .A2(_03112_),
    .B1(_03245_),
    .C1(_03246_),
    .X(_03248_));
 sky130_fd_sc_hd__o211a_1 _09182_ (.A1(_03245_),
    .A2(_03246_),
    .B1(_03065_),
    .C1(_03112_),
    .X(_03249_));
 sky130_fd_sc_hd__a211o_1 _09183_ (.A1(_03107_),
    .A2(_03109_),
    .B1(_03247_),
    .C1(_03249_),
    .X(_03250_));
 sky130_fd_sc_hd__o211ai_2 _09184_ (.A1(_03247_),
    .A2(_03249_),
    .B1(_03107_),
    .C1(_03109_),
    .Y(_03251_));
 sky130_fd_sc_hd__o211ai_2 _09185_ (.A1(_03115_),
    .A2(_03117_),
    .B1(_03250_),
    .C1(_03251_),
    .Y(_03252_));
 sky130_fd_sc_hd__a211o_1 _09186_ (.A1(_03250_),
    .A2(_03251_),
    .B1(_03115_),
    .C1(_03117_),
    .X(_03253_));
 sky130_fd_sc_hd__nand3_1 _09187_ (.A(_03129_),
    .B(_03252_),
    .C(_03253_),
    .Y(_03254_));
 sky130_fd_sc_hd__a21o_1 _09188_ (.A1(_03252_),
    .A2(_03253_),
    .B1(_03129_),
    .X(_03256_));
 sky130_fd_sc_hd__o211a_1 _09189_ (.A1(net129),
    .A2(_03122_),
    .B1(_03254_),
    .C1(_03256_),
    .X(_03257_));
 sky130_fd_sc_hd__a211oi_1 _09190_ (.A1(_03254_),
    .A2(_03256_),
    .B1(net129),
    .C1(_03122_),
    .Y(_03258_));
 sky130_fd_sc_hd__or2_1 _09191_ (.A(_03257_),
    .B(_03258_),
    .X(_03259_));
 sky130_fd_sc_hd__nor2_1 _09192_ (.A(_02989_),
    .B(_03127_),
    .Y(_03260_));
 sky130_fd_sc_hd__nand2_1 _09193_ (.A(_02991_),
    .B(_03260_),
    .Y(_03261_));
 sky130_fd_sc_hd__a21o_1 _09194_ (.A1(_03125_),
    .A2(_03126_),
    .B1(_02987_),
    .X(_03262_));
 sky130_fd_sc_hd__o21a_1 _09195_ (.A1(_03125_),
    .A2(_03126_),
    .B1(_03262_),
    .X(_03263_));
 sky130_fd_sc_hd__nand2_1 _09196_ (.A(_02990_),
    .B(_03260_),
    .Y(_03264_));
 sky130_fd_sc_hd__o211a_2 _09197_ (.A1(_02691_),
    .A2(_03261_),
    .B1(_03263_),
    .C1(_03264_),
    .X(_03265_));
 sky130_fd_sc_hd__a311o_4 _09198_ (.A1(_02041_),
    .A2(_02044_),
    .A3(_02045_),
    .B1(_02692_),
    .C1(_03261_),
    .X(_03267_));
 sky130_fd_sc_hd__a21oi_1 _09199_ (.A1(_03265_),
    .A2(_03267_),
    .B1(_03259_),
    .Y(_03268_));
 sky130_fd_sc_hd__and3_1 _09200_ (.A(_03259_),
    .B(_03265_),
    .C(_03267_),
    .X(_03269_));
 sky130_fd_sc_hd__nor2_1 _09201_ (.A(_03268_),
    .B(_03269_),
    .Y(net99));
 sky130_fd_sc_hd__nor2_1 _09202_ (.A(_03257_),
    .B(_03268_),
    .Y(_03270_));
 sky130_fd_sc_hd__and4_1 _09203_ (.A(net426),
    .B(net422),
    .C(net508),
    .D(net503),
    .X(_03271_));
 sky130_fd_sc_hd__a22oi_1 _09204_ (.A1(net422),
    .A2(net508),
    .B1(net503),
    .B2(net426),
    .Y(_03272_));
 sky130_fd_sc_hd__or2_1 _09205_ (.A(_03271_),
    .B(_03272_),
    .X(_03273_));
 sky130_fd_sc_hd__nand2_1 _09206_ (.A(_03136_),
    .B(_03139_),
    .Y(_03274_));
 sky130_fd_sc_hd__a21o_1 _09207_ (.A1(_03136_),
    .A2(_03139_),
    .B1(_03273_),
    .X(_03275_));
 sky130_fd_sc_hd__xnor2_1 _09208_ (.A(_03273_),
    .B(_03274_),
    .Y(_03277_));
 sky130_fd_sc_hd__and4_1 _09209_ (.A(net412),
    .B(net404),
    .C(net531),
    .D(net522),
    .X(_03278_));
 sky130_fd_sc_hd__a22o_1 _09210_ (.A1(net404),
    .A2(net531),
    .B1(net522),
    .B2(net412),
    .X(_03279_));
 sky130_fd_sc_hd__and2b_1 _09211_ (.A_N(_03278_),
    .B(_03279_),
    .X(_03280_));
 sky130_fd_sc_hd__nand2_1 _09212_ (.A(net397),
    .B(net539),
    .Y(_03281_));
 sky130_fd_sc_hd__xnor2_1 _09213_ (.A(_03280_),
    .B(_03281_),
    .Y(_03282_));
 sky130_fd_sc_hd__nand2_1 _09214_ (.A(_03277_),
    .B(_03282_),
    .Y(_03283_));
 sky130_fd_sc_hd__xor2_1 _09215_ (.A(_03277_),
    .B(_03282_),
    .X(_03284_));
 sky130_fd_sc_hd__o21a_1 _09216_ (.A1(_03141_),
    .A2(_03143_),
    .B1(_03284_),
    .X(_03285_));
 sky130_fd_sc_hd__nor3_1 _09217_ (.A(_03141_),
    .B(_03143_),
    .C(_03284_),
    .Y(_03286_));
 sky130_fd_sc_hd__or2_1 _09218_ (.A(_03285_),
    .B(_03286_),
    .X(_03287_));
 sky130_fd_sc_hd__and4_1 _09219_ (.A(net607),
    .B(net591),
    .C(net327),
    .D(net319),
    .X(_03288_));
 sky130_fd_sc_hd__a22o_1 _09220_ (.A1(net591),
    .A2(net327),
    .B1(net319),
    .B2(net607),
    .X(_03289_));
 sky130_fd_sc_hd__and2b_1 _09221_ (.A_N(_03288_),
    .B(_03289_),
    .X(_03290_));
 sky130_fd_sc_hd__nand2_1 _09222_ (.A(net615),
    .B(net312),
    .Y(_03291_));
 sky130_fd_sc_hd__xnor2_1 _09223_ (.A(_03290_),
    .B(_03291_),
    .Y(_03292_));
 sky130_fd_sc_hd__nand4_1 _09224_ (.A(net357),
    .B(net349),
    .C(net577),
    .D(net571),
    .Y(_03293_));
 sky130_fd_sc_hd__a22o_1 _09225_ (.A1(net349),
    .A2(net577),
    .B1(net571),
    .B2(net357),
    .X(_03294_));
 sky130_fd_sc_hd__and2_1 _09226_ (.A(net335),
    .B(net584),
    .X(_03295_));
 sky130_fd_sc_hd__a21o_1 _09227_ (.A1(_03293_),
    .A2(_03294_),
    .B1(_03295_),
    .X(_03296_));
 sky130_fd_sc_hd__nand3_1 _09228_ (.A(_03293_),
    .B(_03294_),
    .C(_03295_),
    .Y(_03298_));
 sky130_fd_sc_hd__a21bo_1 _09229_ (.A1(_03162_),
    .A2(_03163_),
    .B1_N(_03161_),
    .X(_03299_));
 sky130_fd_sc_hd__and3_1 _09230_ (.A(_03296_),
    .B(_03298_),
    .C(_03299_),
    .X(_03300_));
 sky130_fd_sc_hd__a21o_1 _09231_ (.A1(_03296_),
    .A2(_03298_),
    .B1(_03299_),
    .X(_03301_));
 sky130_fd_sc_hd__and2b_1 _09232_ (.A_N(_03300_),
    .B(_03301_),
    .X(_03302_));
 sky130_fd_sc_hd__xnor2_1 _09233_ (.A(_03292_),
    .B(_03302_),
    .Y(_03303_));
 sky130_fd_sc_hd__nand2_1 _09234_ (.A(_03174_),
    .B(_03177_),
    .Y(_03304_));
 sky130_fd_sc_hd__a31o_1 _09235_ (.A1(net397),
    .A2(net553),
    .A3(_03131_),
    .B1(_03130_),
    .X(_03305_));
 sky130_fd_sc_hd__nand4_1 _09236_ (.A(net389),
    .B(net373),
    .C(net557),
    .D(net553),
    .Y(_03306_));
 sky130_fd_sc_hd__a22o_1 _09237_ (.A1(net373),
    .A2(net557),
    .B1(net553),
    .B2(net389),
    .X(_03307_));
 sky130_fd_sc_hd__a22o_1 _09238_ (.A1(net365),
    .A2(net564),
    .B1(_03306_),
    .B2(_03307_),
    .X(_03309_));
 sky130_fd_sc_hd__nand4_1 _09239_ (.A(net365),
    .B(net564),
    .C(_03306_),
    .D(_03307_),
    .Y(_03310_));
 sky130_fd_sc_hd__nand3_1 _09240_ (.A(_03305_),
    .B(_03309_),
    .C(_03310_),
    .Y(_03311_));
 sky130_fd_sc_hd__a21o_1 _09241_ (.A1(_03309_),
    .A2(_03310_),
    .B1(_03305_),
    .X(_03312_));
 sky130_fd_sc_hd__nand3_1 _09242_ (.A(_03304_),
    .B(_03311_),
    .C(_03312_),
    .Y(_03313_));
 sky130_fd_sc_hd__a21o_1 _09243_ (.A1(_03311_),
    .A2(_03312_),
    .B1(_03304_),
    .X(_03314_));
 sky130_fd_sc_hd__a21bo_1 _09244_ (.A1(_03172_),
    .A2(_03180_),
    .B1_N(_03179_),
    .X(_03315_));
 sky130_fd_sc_hd__and3_1 _09245_ (.A(_03313_),
    .B(_03314_),
    .C(_03315_),
    .X(_03316_));
 sky130_fd_sc_hd__inv_2 _09246_ (.A(_03316_),
    .Y(_03317_));
 sky130_fd_sc_hd__a21oi_1 _09247_ (.A1(_03313_),
    .A2(_03314_),
    .B1(_03315_),
    .Y(_03318_));
 sky130_fd_sc_hd__nor3_1 _09248_ (.A(_03303_),
    .B(_03316_),
    .C(_03318_),
    .Y(_03320_));
 sky130_fd_sc_hd__or3_1 _09249_ (.A(_03303_),
    .B(_03316_),
    .C(_03318_),
    .X(_03321_));
 sky130_fd_sc_hd__o21a_1 _09250_ (.A1(_03316_),
    .A2(_03318_),
    .B1(_03303_),
    .X(_03322_));
 sky130_fd_sc_hd__a211oi_2 _09251_ (.A1(_03147_),
    .A2(_03151_),
    .B1(_03320_),
    .C1(_03322_),
    .Y(_03323_));
 sky130_fd_sc_hd__o211a_1 _09252_ (.A1(_03320_),
    .A2(_03322_),
    .B1(_03147_),
    .C1(_03151_),
    .X(_03324_));
 sky130_fd_sc_hd__a211oi_4 _09253_ (.A1(_03185_),
    .A2(_03188_),
    .B1(_03323_),
    .C1(_03324_),
    .Y(_03325_));
 sky130_fd_sc_hd__o211a_1 _09254_ (.A1(net152),
    .A2(_03324_),
    .B1(_03185_),
    .C1(_03188_),
    .X(_03326_));
 sky130_fd_sc_hd__or3_2 _09255_ (.A(_03287_),
    .B(_03325_),
    .C(_03326_),
    .X(_03327_));
 sky130_fd_sc_hd__o21ai_2 _09256_ (.A1(_03325_),
    .A2(_03326_),
    .B1(_03287_),
    .Y(_03328_));
 sky130_fd_sc_hd__o211ai_4 _09257_ (.A1(_03153_),
    .A2(_03195_),
    .B1(_03327_),
    .C1(_03328_),
    .Y(_03329_));
 sky130_fd_sc_hd__a211o_1 _09258_ (.A1(_03327_),
    .A2(_03328_),
    .B1(_03153_),
    .C1(_03195_),
    .X(_03331_));
 sky130_fd_sc_hd__and4_1 _09259_ (.A(net297),
    .B(net220),
    .C(net276),
    .D(net268),
    .X(_03332_));
 sky130_fd_sc_hd__a22oi_1 _09260_ (.A1(net220),
    .A2(net276),
    .B1(net268),
    .B2(net297),
    .Y(_03333_));
 sky130_fd_sc_hd__o2bb2a_1 _09261_ (.A1_N(net381),
    .A2_N(net260),
    .B1(_03332_),
    .B2(_03333_),
    .X(_03334_));
 sky130_fd_sc_hd__and4bb_1 _09262_ (.A_N(_03332_),
    .B_N(_03333_),
    .C(net381),
    .D(net265),
    .X(_03335_));
 sky130_fd_sc_hd__nor2_1 _09263_ (.A(_03334_),
    .B(_03335_),
    .Y(_03336_));
 sky130_fd_sc_hd__nor2_1 _09264_ (.A(_03201_),
    .B(_03204_),
    .Y(_03337_));
 sky130_fd_sc_hd__and2b_1 _09265_ (.A_N(_03337_),
    .B(_03336_),
    .X(_03338_));
 sky130_fd_sc_hd__xnor2_1 _09266_ (.A(_03336_),
    .B(_03337_),
    .Y(_03339_));
 sky130_fd_sc_hd__and2_1 _09267_ (.A(net464),
    .B(net254),
    .X(_03340_));
 sky130_fd_sc_hd__xnor2_1 _09268_ (.A(_03339_),
    .B(_03340_),
    .Y(_03342_));
 sky130_fd_sc_hd__a21oi_1 _09269_ (.A1(_03208_),
    .A2(_03209_),
    .B1(_03207_),
    .Y(_03343_));
 sky130_fd_sc_hd__xnor2_1 _09270_ (.A(_03342_),
    .B(_03343_),
    .Y(_03344_));
 sky130_fd_sc_hd__nand2_1 _09271_ (.A(net545),
    .B(net246),
    .Y(_03345_));
 sky130_fd_sc_hd__or2_1 _09272_ (.A(_03344_),
    .B(_03345_),
    .X(_03346_));
 sky130_fd_sc_hd__xor2_1 _09273_ (.A(_03344_),
    .B(_03345_),
    .X(_03347_));
 sky130_fd_sc_hd__a21o_1 _09274_ (.A1(_03160_),
    .A2(_03169_),
    .B1(_03168_),
    .X(_03348_));
 sky130_fd_sc_hd__nand2_1 _09275_ (.A(_03221_),
    .B(_03225_),
    .Y(_03349_));
 sky130_fd_sc_hd__a31o_1 _09276_ (.A1(net160),
    .A2(net312),
    .A3(_03157_),
    .B1(_03155_),
    .X(_03350_));
 sky130_fd_sc_hd__nand4_2 _09277_ (.A(net167),
    .B(net160),
    .C(net304),
    .D(net290),
    .Y(_03351_));
 sky130_fd_sc_hd__a22o_1 _09278_ (.A1(net160),
    .A2(net304),
    .B1(net290),
    .B2(net167),
    .X(_03353_));
 sky130_fd_sc_hd__a22o_1 _09279_ (.A1(net175),
    .A2(net283),
    .B1(_03351_),
    .B2(_03353_),
    .X(_03354_));
 sky130_fd_sc_hd__nand4_2 _09280_ (.A(net175),
    .B(net283),
    .C(_03351_),
    .D(_03353_),
    .Y(_03355_));
 sky130_fd_sc_hd__nand3_2 _09281_ (.A(_03350_),
    .B(_03354_),
    .C(_03355_),
    .Y(_03356_));
 sky130_fd_sc_hd__a21o_1 _09282_ (.A1(_03354_),
    .A2(_03355_),
    .B1(_03350_),
    .X(_03357_));
 sky130_fd_sc_hd__nand3_2 _09283_ (.A(_03349_),
    .B(_03356_),
    .C(_03357_),
    .Y(_03358_));
 sky130_fd_sc_hd__a21o_1 _09284_ (.A1(_03356_),
    .A2(_03357_),
    .B1(_03349_),
    .X(_03359_));
 sky130_fd_sc_hd__and3_2 _09285_ (.A(_03348_),
    .B(_03358_),
    .C(_03359_),
    .X(_03360_));
 sky130_fd_sc_hd__a21oi_2 _09286_ (.A1(_03358_),
    .A2(_03359_),
    .B1(_03348_),
    .Y(_03361_));
 sky130_fd_sc_hd__a211oi_4 _09287_ (.A1(_03226_),
    .A2(_03228_),
    .B1(_03360_),
    .C1(_03361_),
    .Y(_03362_));
 sky130_fd_sc_hd__o211a_1 _09288_ (.A1(_03360_),
    .A2(_03361_),
    .B1(_03226_),
    .C1(_03228_),
    .X(_03364_));
 sky130_fd_sc_hd__a211o_1 _09289_ (.A1(_03231_),
    .A2(_03234_),
    .B1(_03362_),
    .C1(_03364_),
    .X(_03365_));
 sky130_fd_sc_hd__inv_2 _09290_ (.A(_03365_),
    .Y(_03366_));
 sky130_fd_sc_hd__o211ai_1 _09291_ (.A1(_03362_),
    .A2(_03364_),
    .B1(_03231_),
    .C1(_03234_),
    .Y(_03367_));
 sky130_fd_sc_hd__and3_1 _09292_ (.A(_03347_),
    .B(_03365_),
    .C(_03367_),
    .X(_03368_));
 sky130_fd_sc_hd__a21oi_1 _09293_ (.A1(_03365_),
    .A2(_03367_),
    .B1(_03347_),
    .Y(_03369_));
 sky130_fd_sc_hd__a211oi_1 _09294_ (.A1(_03191_),
    .A2(_03193_),
    .B1(_03368_),
    .C1(_03369_),
    .Y(_03370_));
 sky130_fd_sc_hd__a211o_1 _09295_ (.A1(_03191_),
    .A2(_03193_),
    .B1(_03368_),
    .C1(_03369_),
    .X(_03371_));
 sky130_fd_sc_hd__o211a_1 _09296_ (.A1(_03368_),
    .A2(_03369_),
    .B1(_03191_),
    .C1(_03193_),
    .X(_03372_));
 sky130_fd_sc_hd__a211o_1 _09297_ (.A1(_03236_),
    .A2(_03238_),
    .B1(_03370_),
    .C1(_03372_),
    .X(_03373_));
 sky130_fd_sc_hd__o211ai_2 _09298_ (.A1(_03370_),
    .A2(_03372_),
    .B1(_03236_),
    .C1(_03238_),
    .Y(_03375_));
 sky130_fd_sc_hd__nand4_2 _09299_ (.A(_03329_),
    .B(_03331_),
    .C(_03373_),
    .D(_03375_),
    .Y(_03376_));
 sky130_fd_sc_hd__a22o_1 _09300_ (.A1(_03329_),
    .A2(_03331_),
    .B1(_03373_),
    .B2(_03375_),
    .X(_03377_));
 sky130_fd_sc_hd__o211a_1 _09301_ (.A1(_03197_),
    .A2(_03245_),
    .B1(_03376_),
    .C1(_03377_),
    .X(_03378_));
 sky130_fd_sc_hd__a211oi_1 _09302_ (.A1(_03376_),
    .A2(_03377_),
    .B1(_03197_),
    .C1(_03245_),
    .Y(_03379_));
 sky130_fd_sc_hd__a211oi_2 _09303_ (.A1(_03240_),
    .A2(_03242_),
    .B1(_03378_),
    .C1(_03379_),
    .Y(_03380_));
 sky130_fd_sc_hd__o211a_1 _09304_ (.A1(_03378_),
    .A2(_03379_),
    .B1(_03240_),
    .C1(_03242_),
    .X(_03381_));
 sky130_fd_sc_hd__a211oi_2 _09305_ (.A1(_03248_),
    .A2(_03250_),
    .B1(_03380_),
    .C1(_03381_),
    .Y(_03382_));
 sky130_fd_sc_hd__inv_2 _09306_ (.A(_03382_),
    .Y(_03383_));
 sky130_fd_sc_hd__o211a_1 _09307_ (.A1(_03380_),
    .A2(_03381_),
    .B1(_03248_),
    .C1(_03250_),
    .X(_03384_));
 sky130_fd_sc_hd__a211oi_1 _09308_ (.A1(_03213_),
    .A2(_03216_),
    .B1(_03382_),
    .C1(_03384_),
    .Y(_03386_));
 sky130_fd_sc_hd__a211o_1 _09309_ (.A1(_03213_),
    .A2(_03216_),
    .B1(_03382_),
    .C1(_03384_),
    .X(_03387_));
 sky130_fd_sc_hd__o211a_1 _09310_ (.A1(_03382_),
    .A2(_03384_),
    .B1(_03213_),
    .C1(_03216_),
    .X(_03388_));
 sky130_fd_sc_hd__a211oi_1 _09311_ (.A1(_03252_),
    .A2(_03254_),
    .B1(_03386_),
    .C1(_03388_),
    .Y(_03389_));
 sky130_fd_sc_hd__o211ai_1 _09312_ (.A1(_03386_),
    .A2(_03388_),
    .B1(_03252_),
    .C1(_03254_),
    .Y(_03390_));
 sky130_fd_sc_hd__and2b_1 _09313_ (.A_N(_03389_),
    .B(_03390_),
    .X(_03391_));
 sky130_fd_sc_hd__inv_2 _09314_ (.A(_03391_),
    .Y(_03392_));
 sky130_fd_sc_hd__xnor2_1 _09315_ (.A(_03270_),
    .B(_03391_),
    .Y(net100));
 sky130_fd_sc_hd__and3_1 _09316_ (.A(net422),
    .B(net503),
    .C(_03001_),
    .X(_03393_));
 sky130_fd_sc_hd__and4_1 _09317_ (.A(net412),
    .B(net404),
    .C(net522),
    .D(net508),
    .X(_03394_));
 sky130_fd_sc_hd__a22o_1 _09318_ (.A1(net404),
    .A2(net522),
    .B1(net508),
    .B2(net412),
    .X(_03396_));
 sky130_fd_sc_hd__and2b_1 _09319_ (.A_N(_03394_),
    .B(_03396_),
    .X(_03397_));
 sky130_fd_sc_hd__nand2_1 _09320_ (.A(net397),
    .B(net531),
    .Y(_03398_));
 sky130_fd_sc_hd__xnor2_1 _09321_ (.A(_03397_),
    .B(_03398_),
    .Y(_03399_));
 sky130_fd_sc_hd__xnor2_1 _09322_ (.A(_03393_),
    .B(_03399_),
    .Y(_03400_));
 sky130_fd_sc_hd__a21oi_2 _09323_ (.A1(_03275_),
    .A2(_03283_),
    .B1(_03400_),
    .Y(_03401_));
 sky130_fd_sc_hd__and3_1 _09324_ (.A(_03275_),
    .B(_03283_),
    .C(_03400_),
    .X(_03402_));
 sky130_fd_sc_hd__or2_1 _09325_ (.A(_03401_),
    .B(_03402_),
    .X(_03403_));
 sky130_fd_sc_hd__and4_1 _09326_ (.A(net591),
    .B(net584),
    .C(net327),
    .D(net319),
    .X(_03404_));
 sky130_fd_sc_hd__a22o_1 _09327_ (.A1(net584),
    .A2(net327),
    .B1(net319),
    .B2(net591),
    .X(_03405_));
 sky130_fd_sc_hd__and2b_1 _09328_ (.A_N(_03404_),
    .B(_03405_),
    .X(_03407_));
 sky130_fd_sc_hd__nand2_1 _09329_ (.A(net607),
    .B(net312),
    .Y(_03408_));
 sky130_fd_sc_hd__xnor2_1 _09330_ (.A(_03407_),
    .B(_03408_),
    .Y(_03409_));
 sky130_fd_sc_hd__nand4_1 _09331_ (.A(net357),
    .B(net349),
    .C(net571),
    .D(net564),
    .Y(_03410_));
 sky130_fd_sc_hd__a22o_1 _09332_ (.A1(net349),
    .A2(net571),
    .B1(net564),
    .B2(net357),
    .X(_03411_));
 sky130_fd_sc_hd__and2_1 _09333_ (.A(net335),
    .B(net577),
    .X(_03412_));
 sky130_fd_sc_hd__a21o_1 _09334_ (.A1(_03410_),
    .A2(_03411_),
    .B1(_03412_),
    .X(_03413_));
 sky130_fd_sc_hd__nand3_1 _09335_ (.A(_03410_),
    .B(_03411_),
    .C(_03412_),
    .Y(_03414_));
 sky130_fd_sc_hd__a21bo_1 _09336_ (.A1(_03294_),
    .A2(_03295_),
    .B1_N(_03293_),
    .X(_03415_));
 sky130_fd_sc_hd__and3_1 _09337_ (.A(_03413_),
    .B(_03414_),
    .C(_03415_),
    .X(_03416_));
 sky130_fd_sc_hd__a21o_1 _09338_ (.A1(_03413_),
    .A2(_03414_),
    .B1(_03415_),
    .X(_03418_));
 sky130_fd_sc_hd__and2b_1 _09339_ (.A_N(_03416_),
    .B(_03418_),
    .X(_03419_));
 sky130_fd_sc_hd__xnor2_1 _09340_ (.A(_03409_),
    .B(_03419_),
    .Y(_03420_));
 sky130_fd_sc_hd__nand2_1 _09341_ (.A(_03306_),
    .B(_03310_),
    .Y(_03421_));
 sky130_fd_sc_hd__a31o_1 _09342_ (.A1(net397),
    .A2(net539),
    .A3(_03279_),
    .B1(_03278_),
    .X(_03422_));
 sky130_fd_sc_hd__nand4_1 _09343_ (.A(net389),
    .B(net373),
    .C(net550),
    .D(net536),
    .Y(_03423_));
 sky130_fd_sc_hd__a22o_1 _09344_ (.A1(net373),
    .A2(net550),
    .B1(net536),
    .B2(net389),
    .X(_03424_));
 sky130_fd_sc_hd__a22o_1 _09345_ (.A1(net365),
    .A2(net557),
    .B1(_03423_),
    .B2(_03424_),
    .X(_03425_));
 sky130_fd_sc_hd__nand4_1 _09346_ (.A(net365),
    .B(net557),
    .C(_03423_),
    .D(_03424_),
    .Y(_03426_));
 sky130_fd_sc_hd__nand3_1 _09347_ (.A(_03422_),
    .B(_03425_),
    .C(_03426_),
    .Y(_03427_));
 sky130_fd_sc_hd__a21o_1 _09348_ (.A1(_03425_),
    .A2(_03426_),
    .B1(_03422_),
    .X(_03429_));
 sky130_fd_sc_hd__nand3_1 _09349_ (.A(_03421_),
    .B(_03427_),
    .C(_03429_),
    .Y(_03430_));
 sky130_fd_sc_hd__a21o_1 _09350_ (.A1(_03427_),
    .A2(_03429_),
    .B1(_03421_),
    .X(_03431_));
 sky130_fd_sc_hd__a21bo_1 _09351_ (.A1(_03304_),
    .A2(_03312_),
    .B1_N(_03311_),
    .X(_03432_));
 sky130_fd_sc_hd__and3_1 _09352_ (.A(_03430_),
    .B(_03431_),
    .C(_03432_),
    .X(_03433_));
 sky130_fd_sc_hd__nand3_1 _09353_ (.A(_03430_),
    .B(_03431_),
    .C(_03432_),
    .Y(_03434_));
 sky130_fd_sc_hd__a21oi_1 _09354_ (.A1(_03430_),
    .A2(_03431_),
    .B1(_03432_),
    .Y(_03435_));
 sky130_fd_sc_hd__or3_1 _09355_ (.A(_03420_),
    .B(_03433_),
    .C(_03435_),
    .X(_03436_));
 sky130_fd_sc_hd__o21ai_1 _09356_ (.A1(_03433_),
    .A2(_03435_),
    .B1(_03420_),
    .Y(_03437_));
 sky130_fd_sc_hd__and3_2 _09357_ (.A(_03285_),
    .B(_03436_),
    .C(_03437_),
    .X(_03438_));
 sky130_fd_sc_hd__a21oi_1 _09358_ (.A1(_03436_),
    .A2(_03437_),
    .B1(_03285_),
    .Y(_03440_));
 sky130_fd_sc_hd__a211oi_2 _09359_ (.A1(_03317_),
    .A2(_03321_),
    .B1(_03438_),
    .C1(_03440_),
    .Y(_03441_));
 sky130_fd_sc_hd__o211a_1 _09360_ (.A1(_03438_),
    .A2(_03440_),
    .B1(_03317_),
    .C1(_03321_),
    .X(_03442_));
 sky130_fd_sc_hd__nor3_1 _09361_ (.A(_03403_),
    .B(_03441_),
    .C(_03442_),
    .Y(_03443_));
 sky130_fd_sc_hd__o21a_1 _09362_ (.A1(_03441_),
    .A2(_03442_),
    .B1(_03403_),
    .X(_03444_));
 sky130_fd_sc_hd__o21a_1 _09363_ (.A1(_03443_),
    .A2(_03444_),
    .B1(_03327_),
    .X(_03445_));
 sky130_fd_sc_hd__nor3_1 _09364_ (.A(_03327_),
    .B(_03443_),
    .C(_03444_),
    .Y(_03446_));
 sky130_fd_sc_hd__and4_1 _09365_ (.A(net220),
    .B(net175),
    .C(net275),
    .D(net266),
    .X(_03447_));
 sky130_fd_sc_hd__a22oi_1 _09366_ (.A1(net175),
    .A2(net275),
    .B1(net266),
    .B2(net220),
    .Y(_03448_));
 sky130_fd_sc_hd__o2bb2a_1 _09367_ (.A1_N(net297),
    .A2_N(net259),
    .B1(_03447_),
    .B2(_03448_),
    .X(_03449_));
 sky130_fd_sc_hd__and4bb_1 _09368_ (.A_N(_03447_),
    .B_N(_03448_),
    .C(net297),
    .D(net259),
    .X(_03451_));
 sky130_fd_sc_hd__nor2_1 _09369_ (.A(_03449_),
    .B(_03451_),
    .Y(_03452_));
 sky130_fd_sc_hd__nor2_1 _09370_ (.A(_03332_),
    .B(_03335_),
    .Y(_03453_));
 sky130_fd_sc_hd__and2b_1 _09371_ (.A_N(_03453_),
    .B(_03452_),
    .X(_03454_));
 sky130_fd_sc_hd__xnor2_1 _09372_ (.A(_03452_),
    .B(_03453_),
    .Y(_03455_));
 sky130_fd_sc_hd__and2_1 _09373_ (.A(net381),
    .B(net254),
    .X(_03456_));
 sky130_fd_sc_hd__xnor2_1 _09374_ (.A(_03455_),
    .B(_03456_),
    .Y(_03457_));
 sky130_fd_sc_hd__a21oi_1 _09375_ (.A1(_03339_),
    .A2(_03340_),
    .B1(_03338_),
    .Y(_03458_));
 sky130_fd_sc_hd__or2_1 _09376_ (.A(_03457_),
    .B(_03458_),
    .X(_03459_));
 sky130_fd_sc_hd__xnor2_1 _09377_ (.A(_03457_),
    .B(_03458_),
    .Y(_03460_));
 sky130_fd_sc_hd__nand2_1 _09378_ (.A(net464),
    .B(net246),
    .Y(_03462_));
 sky130_fd_sc_hd__or2_1 _09379_ (.A(_03460_),
    .B(_03462_),
    .X(_03463_));
 sky130_fd_sc_hd__xor2_1 _09380_ (.A(_03460_),
    .B(_03462_),
    .X(_03464_));
 sky130_fd_sc_hd__a21o_1 _09381_ (.A1(_03292_),
    .A2(_03301_),
    .B1(_03300_),
    .X(_03465_));
 sky130_fd_sc_hd__nand2_1 _09382_ (.A(_03351_),
    .B(_03355_),
    .Y(_03466_));
 sky130_fd_sc_hd__a31o_1 _09383_ (.A1(net615),
    .A2(net312),
    .A3(_03289_),
    .B1(_03288_),
    .X(_03467_));
 sky130_fd_sc_hd__nand4_2 _09384_ (.A(net159),
    .B(net615),
    .C(net304),
    .D(net290),
    .Y(_03468_));
 sky130_fd_sc_hd__a22o_1 _09385_ (.A1(net615),
    .A2(net304),
    .B1(net290),
    .B2(net159),
    .X(_03469_));
 sky130_fd_sc_hd__a22o_1 _09386_ (.A1(net167),
    .A2(net283),
    .B1(_03468_),
    .B2(_03469_),
    .X(_03470_));
 sky130_fd_sc_hd__nand4_2 _09387_ (.A(net167),
    .B(net283),
    .C(_03468_),
    .D(_03469_),
    .Y(_03471_));
 sky130_fd_sc_hd__nand3_2 _09388_ (.A(_03467_),
    .B(_03470_),
    .C(_03471_),
    .Y(_03473_));
 sky130_fd_sc_hd__a21o_1 _09389_ (.A1(_03470_),
    .A2(_03471_),
    .B1(_03467_),
    .X(_03474_));
 sky130_fd_sc_hd__nand3_2 _09390_ (.A(_03466_),
    .B(_03473_),
    .C(_03474_),
    .Y(_03475_));
 sky130_fd_sc_hd__a21o_1 _09391_ (.A1(_03473_),
    .A2(_03474_),
    .B1(_03466_),
    .X(_03476_));
 sky130_fd_sc_hd__and3_1 _09392_ (.A(_03465_),
    .B(_03475_),
    .C(_03476_),
    .X(_03477_));
 sky130_fd_sc_hd__nand3_1 _09393_ (.A(_03465_),
    .B(_03475_),
    .C(_03476_),
    .Y(_03478_));
 sky130_fd_sc_hd__a21oi_1 _09394_ (.A1(_03475_),
    .A2(_03476_),
    .B1(_03465_),
    .Y(_03479_));
 sky130_fd_sc_hd__a211o_2 _09395_ (.A1(_03356_),
    .A2(_03358_),
    .B1(_03477_),
    .C1(_03479_),
    .X(_03480_));
 sky130_fd_sc_hd__o211ai_2 _09396_ (.A1(_03477_),
    .A2(_03479_),
    .B1(_03356_),
    .C1(_03358_),
    .Y(_03481_));
 sky130_fd_sc_hd__o211ai_4 _09397_ (.A1(_03360_),
    .A2(_03362_),
    .B1(_03480_),
    .C1(_03481_),
    .Y(_03482_));
 sky130_fd_sc_hd__a211o_1 _09398_ (.A1(_03480_),
    .A2(_03481_),
    .B1(_03360_),
    .C1(_03362_),
    .X(_03484_));
 sky130_fd_sc_hd__nand3_2 _09399_ (.A(_03464_),
    .B(_03482_),
    .C(_03484_),
    .Y(_03485_));
 sky130_fd_sc_hd__a21o_1 _09400_ (.A1(_03482_),
    .A2(_03484_),
    .B1(_03464_),
    .X(_03486_));
 sky130_fd_sc_hd__o211ai_4 _09401_ (.A1(net152),
    .A2(_03325_),
    .B1(_03485_),
    .C1(_03486_),
    .Y(_03487_));
 sky130_fd_sc_hd__a211o_1 _09402_ (.A1(_03485_),
    .A2(_03486_),
    .B1(net152),
    .C1(_03325_),
    .X(_03488_));
 sky130_fd_sc_hd__o211ai_2 _09403_ (.A1(_03366_),
    .A2(_03368_),
    .B1(_03487_),
    .C1(_03488_),
    .Y(_03489_));
 sky130_fd_sc_hd__a211o_1 _09404_ (.A1(_03487_),
    .A2(_03488_),
    .B1(_03366_),
    .C1(_03368_),
    .X(_03490_));
 sky130_fd_sc_hd__and4bb_1 _09405_ (.A_N(_03445_),
    .B_N(_03446_),
    .C(_03489_),
    .D(_03490_),
    .X(_03491_));
 sky130_fd_sc_hd__a2bb2oi_1 _09406_ (.A1_N(_03445_),
    .A2_N(_03446_),
    .B1(_03489_),
    .B2(_03490_),
    .Y(_03492_));
 sky130_fd_sc_hd__a211oi_2 _09407_ (.A1(_03329_),
    .A2(_03376_),
    .B1(_03491_),
    .C1(_03492_),
    .Y(_03493_));
 sky130_fd_sc_hd__inv_2 _09408_ (.A(_03493_),
    .Y(_03495_));
 sky130_fd_sc_hd__o211a_1 _09409_ (.A1(_03491_),
    .A2(_03492_),
    .B1(_03329_),
    .C1(_03376_),
    .X(_03496_));
 sky130_fd_sc_hd__a211o_1 _09410_ (.A1(_03371_),
    .A2(_03373_),
    .B1(_03493_),
    .C1(_03496_),
    .X(_03497_));
 sky130_fd_sc_hd__o211ai_2 _09411_ (.A1(_03493_),
    .A2(_03496_),
    .B1(_03371_),
    .C1(_03373_),
    .Y(_03498_));
 sky130_fd_sc_hd__o211ai_2 _09412_ (.A1(_03378_),
    .A2(_03380_),
    .B1(_03497_),
    .C1(_03498_),
    .Y(_03499_));
 sky130_fd_sc_hd__a211o_1 _09413_ (.A1(_03497_),
    .A2(_03498_),
    .B1(_03378_),
    .C1(_03380_),
    .X(_03500_));
 sky130_fd_sc_hd__o21ai_1 _09414_ (.A1(_03342_),
    .A2(_03343_),
    .B1(_03346_),
    .Y(_03501_));
 sky130_fd_sc_hd__and3_1 _09415_ (.A(_03499_),
    .B(_03500_),
    .C(_03501_),
    .X(_03502_));
 sky130_fd_sc_hd__nand3_1 _09416_ (.A(_03499_),
    .B(_03500_),
    .C(_03501_),
    .Y(_03503_));
 sky130_fd_sc_hd__a21oi_1 _09417_ (.A1(_03499_),
    .A2(_03500_),
    .B1(_03501_),
    .Y(_03504_));
 sky130_fd_sc_hd__a211oi_2 _09418_ (.A1(_03383_),
    .A2(_03387_),
    .B1(_03502_),
    .C1(_03504_),
    .Y(_03506_));
 sky130_fd_sc_hd__o211a_1 _09419_ (.A1(_03502_),
    .A2(_03504_),
    .B1(_03383_),
    .C1(_03387_),
    .X(_03507_));
 sky130_fd_sc_hd__nor2_1 _09420_ (.A(_03506_),
    .B(_03507_),
    .Y(_03508_));
 sky130_fd_sc_hd__o21a_1 _09421_ (.A1(_03257_),
    .A2(_03389_),
    .B1(_03390_),
    .X(_03509_));
 sky130_fd_sc_hd__a21o_1 _09422_ (.A1(_03268_),
    .A2(_03391_),
    .B1(_03509_),
    .X(_03510_));
 sky130_fd_sc_hd__xor2_1 _09423_ (.A(_03508_),
    .B(_03510_),
    .X(net101));
 sky130_fd_sc_hd__and4_1 _09424_ (.A(net412),
    .B(net404),
    .C(net508),
    .D(net503),
    .X(_03511_));
 sky130_fd_sc_hd__a22o_1 _09425_ (.A1(net404),
    .A2(net508),
    .B1(net503),
    .B2(net412),
    .X(_03512_));
 sky130_fd_sc_hd__and2b_1 _09426_ (.A_N(_03511_),
    .B(_03512_),
    .X(_03513_));
 sky130_fd_sc_hd__nand2_1 _09427_ (.A(net397),
    .B(net521),
    .Y(_03514_));
 sky130_fd_sc_hd__xnor2_1 _09428_ (.A(_03513_),
    .B(_03514_),
    .Y(_03516_));
 sky130_fd_sc_hd__a21oi_1 _09429_ (.A1(_03393_),
    .A2(_03399_),
    .B1(_03271_),
    .Y(_03517_));
 sky130_fd_sc_hd__and2b_1 _09430_ (.A_N(_03517_),
    .B(_03516_),
    .X(_03518_));
 sky130_fd_sc_hd__and2b_1 _09431_ (.A_N(_03516_),
    .B(_03517_),
    .X(_03519_));
 sky130_fd_sc_hd__nor2_1 _09432_ (.A(_03518_),
    .B(_03519_),
    .Y(_03520_));
 sky130_fd_sc_hd__and4_1 _09433_ (.A(net584),
    .B(net327),
    .C(net577),
    .D(net319),
    .X(_03521_));
 sky130_fd_sc_hd__a22o_1 _09434_ (.A1(net327),
    .A2(net577),
    .B1(net319),
    .B2(net584),
    .X(_03522_));
 sky130_fd_sc_hd__and2b_1 _09435_ (.A_N(_03521_),
    .B(_03522_),
    .X(_03523_));
 sky130_fd_sc_hd__nand2_1 _09436_ (.A(net591),
    .B(net312),
    .Y(_03524_));
 sky130_fd_sc_hd__xnor2_1 _09437_ (.A(_03523_),
    .B(_03524_),
    .Y(_03525_));
 sky130_fd_sc_hd__nand4_1 _09438_ (.A(net357),
    .B(net349),
    .C(net564),
    .D(net557),
    .Y(_03527_));
 sky130_fd_sc_hd__a22o_1 _09439_ (.A1(net349),
    .A2(net564),
    .B1(net557),
    .B2(net357),
    .X(_03528_));
 sky130_fd_sc_hd__and2_1 _09440_ (.A(net335),
    .B(net571),
    .X(_03529_));
 sky130_fd_sc_hd__a21o_1 _09441_ (.A1(_03527_),
    .A2(_03528_),
    .B1(_03529_),
    .X(_03530_));
 sky130_fd_sc_hd__nand3_1 _09442_ (.A(_03527_),
    .B(_03528_),
    .C(_03529_),
    .Y(_03531_));
 sky130_fd_sc_hd__a21bo_1 _09443_ (.A1(_03411_),
    .A2(_03412_),
    .B1_N(_03410_),
    .X(_03532_));
 sky130_fd_sc_hd__and3_1 _09444_ (.A(_03530_),
    .B(_03531_),
    .C(_03532_),
    .X(_03533_));
 sky130_fd_sc_hd__a21o_1 _09445_ (.A1(_03530_),
    .A2(_03531_),
    .B1(_03532_),
    .X(_03534_));
 sky130_fd_sc_hd__and2b_1 _09446_ (.A_N(_03533_),
    .B(_03534_),
    .X(_03535_));
 sky130_fd_sc_hd__xnor2_1 _09447_ (.A(_03525_),
    .B(_03535_),
    .Y(_03536_));
 sky130_fd_sc_hd__nand2_1 _09448_ (.A(_03423_),
    .B(_03426_),
    .Y(_03538_));
 sky130_fd_sc_hd__a31o_1 _09449_ (.A1(net397),
    .A2(net531),
    .A3(_03396_),
    .B1(_03394_),
    .X(_03539_));
 sky130_fd_sc_hd__nand4_1 _09450_ (.A(net389),
    .B(net373),
    .C(net536),
    .D(net529),
    .Y(_03540_));
 sky130_fd_sc_hd__a22o_1 _09451_ (.A1(net373),
    .A2(net536),
    .B1(net529),
    .B2(net389),
    .X(_03541_));
 sky130_fd_sc_hd__a22o_1 _09452_ (.A1(net365),
    .A2(net550),
    .B1(_03540_),
    .B2(_03541_),
    .X(_03542_));
 sky130_fd_sc_hd__nand4_1 _09453_ (.A(net365),
    .B(net550),
    .C(_03540_),
    .D(_03541_),
    .Y(_03543_));
 sky130_fd_sc_hd__nand3_1 _09454_ (.A(_03539_),
    .B(_03542_),
    .C(_03543_),
    .Y(_03544_));
 sky130_fd_sc_hd__a21o_1 _09455_ (.A1(_03542_),
    .A2(_03543_),
    .B1(_03539_),
    .X(_03545_));
 sky130_fd_sc_hd__nand3_1 _09456_ (.A(_03538_),
    .B(_03544_),
    .C(_03545_),
    .Y(_03546_));
 sky130_fd_sc_hd__a21o_1 _09457_ (.A1(_03544_),
    .A2(_03545_),
    .B1(_03538_),
    .X(_03547_));
 sky130_fd_sc_hd__a21bo_1 _09458_ (.A1(_03421_),
    .A2(_03429_),
    .B1_N(_03427_),
    .X(_03549_));
 sky130_fd_sc_hd__and3_1 _09459_ (.A(_03546_),
    .B(_03547_),
    .C(_03549_),
    .X(_03550_));
 sky130_fd_sc_hd__nand3_1 _09460_ (.A(_03546_),
    .B(_03547_),
    .C(_03549_),
    .Y(_03551_));
 sky130_fd_sc_hd__a21oi_1 _09461_ (.A1(_03546_),
    .A2(_03547_),
    .B1(_03549_),
    .Y(_03552_));
 sky130_fd_sc_hd__or3_2 _09462_ (.A(_03536_),
    .B(_03550_),
    .C(_03552_),
    .X(_03553_));
 sky130_fd_sc_hd__o21ai_1 _09463_ (.A1(_03550_),
    .A2(_03552_),
    .B1(_03536_),
    .Y(_03554_));
 sky130_fd_sc_hd__and3_1 _09464_ (.A(_03401_),
    .B(_03553_),
    .C(_03554_),
    .X(_03555_));
 sky130_fd_sc_hd__nand3_1 _09465_ (.A(_03401_),
    .B(_03553_),
    .C(_03554_),
    .Y(_03556_));
 sky130_fd_sc_hd__a21oi_1 _09466_ (.A1(_03553_),
    .A2(_03554_),
    .B1(_03401_),
    .Y(_03557_));
 sky130_fd_sc_hd__a211o_1 _09467_ (.A1(_03434_),
    .A2(_03436_),
    .B1(_03555_),
    .C1(_03557_),
    .X(_03558_));
 sky130_fd_sc_hd__o211ai_1 _09468_ (.A1(_03555_),
    .A2(_03557_),
    .B1(_03434_),
    .C1(_03436_),
    .Y(_03560_));
 sky130_fd_sc_hd__and3_1 _09469_ (.A(_03520_),
    .B(_03558_),
    .C(_03560_),
    .X(_03561_));
 sky130_fd_sc_hd__a21oi_1 _09470_ (.A1(_03558_),
    .A2(_03560_),
    .B1(_03520_),
    .Y(_03562_));
 sky130_fd_sc_hd__o21bai_1 _09471_ (.A1(_03561_),
    .A2(_03562_),
    .B1_N(_03443_),
    .Y(_03563_));
 sky130_fd_sc_hd__or3b_2 _09472_ (.A(_03561_),
    .B(_03562_),
    .C_N(_03443_),
    .X(_03564_));
 sky130_fd_sc_hd__and4_1 _09473_ (.A(net175),
    .B(net167),
    .C(net275),
    .D(net266),
    .X(_03565_));
 sky130_fd_sc_hd__a22oi_1 _09474_ (.A1(net167),
    .A2(net275),
    .B1(net266),
    .B2(net175),
    .Y(_03566_));
 sky130_fd_sc_hd__o2bb2a_1 _09475_ (.A1_N(net220),
    .A2_N(net259),
    .B1(_03565_),
    .B2(_03566_),
    .X(_03567_));
 sky130_fd_sc_hd__and4bb_1 _09476_ (.A_N(_03565_),
    .B_N(_03566_),
    .C(net220),
    .D(net259),
    .X(_03568_));
 sky130_fd_sc_hd__nor2_1 _09477_ (.A(_03567_),
    .B(_03568_),
    .Y(_03569_));
 sky130_fd_sc_hd__nor2_1 _09478_ (.A(_03447_),
    .B(_03451_),
    .Y(_03571_));
 sky130_fd_sc_hd__and2b_1 _09479_ (.A_N(_03571_),
    .B(_03569_),
    .X(_03572_));
 sky130_fd_sc_hd__xnor2_1 _09480_ (.A(_03569_),
    .B(_03571_),
    .Y(_03573_));
 sky130_fd_sc_hd__and2_1 _09481_ (.A(net297),
    .B(net249),
    .X(_03574_));
 sky130_fd_sc_hd__xnor2_1 _09482_ (.A(_03573_),
    .B(_03574_),
    .Y(_03575_));
 sky130_fd_sc_hd__a21oi_1 _09483_ (.A1(_03455_),
    .A2(_03456_),
    .B1(_03454_),
    .Y(_03576_));
 sky130_fd_sc_hd__xnor2_1 _09484_ (.A(_03575_),
    .B(_03576_),
    .Y(_03577_));
 sky130_fd_sc_hd__nand2_1 _09485_ (.A(net381),
    .B(net246),
    .Y(_03578_));
 sky130_fd_sc_hd__or2_1 _09486_ (.A(_03577_),
    .B(_03578_),
    .X(_03579_));
 sky130_fd_sc_hd__xor2_1 _09487_ (.A(_03577_),
    .B(_03578_),
    .X(_03580_));
 sky130_fd_sc_hd__a21o_1 _09488_ (.A1(_03409_),
    .A2(_03418_),
    .B1(_03416_),
    .X(_03582_));
 sky130_fd_sc_hd__nand2_1 _09489_ (.A(_03468_),
    .B(_03471_),
    .Y(_03583_));
 sky130_fd_sc_hd__a31o_1 _09490_ (.A1(net607),
    .A2(net312),
    .A3(_03405_),
    .B1(_03404_),
    .X(_03584_));
 sky130_fd_sc_hd__nand4_2 _09491_ (.A(net615),
    .B(net607),
    .C(net304),
    .D(net290),
    .Y(_03585_));
 sky130_fd_sc_hd__a22o_1 _09492_ (.A1(net607),
    .A2(net304),
    .B1(net290),
    .B2(net615),
    .X(_03586_));
 sky130_fd_sc_hd__a22o_1 _09493_ (.A1(net159),
    .A2(net283),
    .B1(_03585_),
    .B2(_03586_),
    .X(_03587_));
 sky130_fd_sc_hd__nand4_2 _09494_ (.A(net159),
    .B(net283),
    .C(_03585_),
    .D(_03586_),
    .Y(_03588_));
 sky130_fd_sc_hd__nand3_2 _09495_ (.A(_03584_),
    .B(_03587_),
    .C(_03588_),
    .Y(_03589_));
 sky130_fd_sc_hd__a21o_1 _09496_ (.A1(_03587_),
    .A2(_03588_),
    .B1(_03584_),
    .X(_03590_));
 sky130_fd_sc_hd__nand3_1 _09497_ (.A(_03583_),
    .B(_03589_),
    .C(_03590_),
    .Y(_03591_));
 sky130_fd_sc_hd__a21o_1 _09498_ (.A1(_03589_),
    .A2(_03590_),
    .B1(_03583_),
    .X(_03593_));
 sky130_fd_sc_hd__and3_1 _09499_ (.A(_03582_),
    .B(_03591_),
    .C(_03593_),
    .X(_03594_));
 sky130_fd_sc_hd__a21oi_1 _09500_ (.A1(_03591_),
    .A2(_03593_),
    .B1(_03582_),
    .Y(_03595_));
 sky130_fd_sc_hd__a211oi_2 _09501_ (.A1(_03473_),
    .A2(_03475_),
    .B1(_03594_),
    .C1(_03595_),
    .Y(_03596_));
 sky130_fd_sc_hd__o211a_1 _09502_ (.A1(_03594_),
    .A2(_03595_),
    .B1(_03473_),
    .C1(_03475_),
    .X(_03597_));
 sky130_fd_sc_hd__a211o_1 _09503_ (.A1(_03478_),
    .A2(_03480_),
    .B1(_03596_),
    .C1(_03597_),
    .X(_03598_));
 sky130_fd_sc_hd__o211ai_1 _09504_ (.A1(_03596_),
    .A2(_03597_),
    .B1(_03478_),
    .C1(_03480_),
    .Y(_03599_));
 sky130_fd_sc_hd__nand3_1 _09505_ (.A(_03580_),
    .B(_03598_),
    .C(_03599_),
    .Y(_03600_));
 sky130_fd_sc_hd__a21o_1 _09506_ (.A1(_03598_),
    .A2(_03599_),
    .B1(_03580_),
    .X(_03601_));
 sky130_fd_sc_hd__o211a_1 _09507_ (.A1(_03438_),
    .A2(_03441_),
    .B1(_03600_),
    .C1(_03601_),
    .X(_03602_));
 sky130_fd_sc_hd__o211ai_1 _09508_ (.A1(_03438_),
    .A2(_03441_),
    .B1(_03600_),
    .C1(_03601_),
    .Y(_03604_));
 sky130_fd_sc_hd__a211oi_1 _09509_ (.A1(_03600_),
    .A2(_03601_),
    .B1(_03438_),
    .C1(_03441_),
    .Y(_03605_));
 sky130_fd_sc_hd__a211o_1 _09510_ (.A1(_03482_),
    .A2(_03485_),
    .B1(_03602_),
    .C1(_03605_),
    .X(_03606_));
 sky130_fd_sc_hd__o211ai_2 _09511_ (.A1(_03602_),
    .A2(_03605_),
    .B1(_03482_),
    .C1(_03485_),
    .Y(_03607_));
 sky130_fd_sc_hd__nand4_2 _09512_ (.A(_03563_),
    .B(_03564_),
    .C(_03606_),
    .D(_03607_),
    .Y(_03608_));
 sky130_fd_sc_hd__a22o_1 _09513_ (.A1(_03563_),
    .A2(_03564_),
    .B1(_03606_),
    .B2(_03607_),
    .X(_03609_));
 sky130_fd_sc_hd__o211a_1 _09514_ (.A1(_03446_),
    .A2(_03491_),
    .B1(_03608_),
    .C1(_03609_),
    .X(_03610_));
 sky130_fd_sc_hd__a211oi_1 _09515_ (.A1(_03608_),
    .A2(_03609_),
    .B1(_03446_),
    .C1(_03491_),
    .Y(_03611_));
 sky130_fd_sc_hd__a211oi_2 _09516_ (.A1(_03487_),
    .A2(_03489_),
    .B1(_03610_),
    .C1(_03611_),
    .Y(_03612_));
 sky130_fd_sc_hd__o211a_1 _09517_ (.A1(_03610_),
    .A2(_03611_),
    .B1(_03487_),
    .C1(_03489_),
    .X(_03613_));
 sky130_fd_sc_hd__a211oi_2 _09518_ (.A1(_03495_),
    .A2(_03497_),
    .B1(_03612_),
    .C1(_03613_),
    .Y(_03615_));
 sky130_fd_sc_hd__o211a_1 _09519_ (.A1(_03612_),
    .A2(_03613_),
    .B1(_03495_),
    .C1(_03497_),
    .X(_03616_));
 sky130_fd_sc_hd__a211oi_2 _09520_ (.A1(_03459_),
    .A2(_03463_),
    .B1(_03615_),
    .C1(_03616_),
    .Y(_03617_));
 sky130_fd_sc_hd__o211a_1 _09521_ (.A1(_03615_),
    .A2(_03616_),
    .B1(_03459_),
    .C1(_03463_),
    .X(_03618_));
 sky130_fd_sc_hd__o211a_1 _09522_ (.A1(_03617_),
    .A2(_03618_),
    .B1(_03499_),
    .C1(_03503_),
    .X(_03619_));
 sky130_fd_sc_hd__a211oi_1 _09523_ (.A1(_03499_),
    .A2(_03503_),
    .B1(_03617_),
    .C1(_03618_),
    .Y(_03620_));
 sky130_fd_sc_hd__nor2_1 _09524_ (.A(_03619_),
    .B(_03620_),
    .Y(_03621_));
 sky130_fd_sc_hd__a21oi_1 _09525_ (.A1(_03508_),
    .A2(_03510_),
    .B1(_03506_),
    .Y(_03622_));
 sky130_fd_sc_hd__xnor2_1 _09526_ (.A(_03621_),
    .B(_03622_),
    .Y(net102));
 sky130_fd_sc_hd__a22o_1 _09527_ (.A1(net397),
    .A2(net507),
    .B1(net501),
    .B2(net404),
    .X(_03623_));
 sky130_fd_sc_hd__nand2_1 _09528_ (.A(net397),
    .B(net501),
    .Y(_03625_));
 sky130_fd_sc_hd__nand4_2 _09529_ (.A(net405),
    .B(net397),
    .C(net508),
    .D(net503),
    .Y(_03626_));
 sky130_fd_sc_hd__and4_1 _09530_ (.A(net327),
    .B(net577),
    .C(net319),
    .D(net571),
    .X(_03627_));
 sky130_fd_sc_hd__a22o_1 _09531_ (.A1(net577),
    .A2(net319),
    .B1(net571),
    .B2(net327),
    .X(_03628_));
 sky130_fd_sc_hd__and2b_1 _09532_ (.A_N(_03627_),
    .B(_03628_),
    .X(_03629_));
 sky130_fd_sc_hd__nand2_1 _09533_ (.A(net584),
    .B(net312),
    .Y(_03630_));
 sky130_fd_sc_hd__xnor2_1 _09534_ (.A(_03629_),
    .B(_03630_),
    .Y(_03631_));
 sky130_fd_sc_hd__nand4_1 _09535_ (.A(net358),
    .B(net350),
    .C(net557),
    .D(net550),
    .Y(_03632_));
 sky130_fd_sc_hd__a22o_1 _09536_ (.A1(net350),
    .A2(net557),
    .B1(net550),
    .B2(net358),
    .X(_03633_));
 sky130_fd_sc_hd__and2_1 _09537_ (.A(net335),
    .B(net564),
    .X(_03634_));
 sky130_fd_sc_hd__a21o_1 _09538_ (.A1(_03632_),
    .A2(_03633_),
    .B1(_03634_),
    .X(_03636_));
 sky130_fd_sc_hd__nand3_1 _09539_ (.A(_03632_),
    .B(_03633_),
    .C(_03634_),
    .Y(_03637_));
 sky130_fd_sc_hd__a21bo_1 _09540_ (.A1(_03528_),
    .A2(_03529_),
    .B1_N(_03527_),
    .X(_03638_));
 sky130_fd_sc_hd__and3_1 _09541_ (.A(_03636_),
    .B(_03637_),
    .C(_03638_),
    .X(_03639_));
 sky130_fd_sc_hd__a21o_1 _09542_ (.A1(_03636_),
    .A2(_03637_),
    .B1(_03638_),
    .X(_03640_));
 sky130_fd_sc_hd__and2b_1 _09543_ (.A_N(_03639_),
    .B(_03640_),
    .X(_03641_));
 sky130_fd_sc_hd__xnor2_1 _09544_ (.A(_03631_),
    .B(_03641_),
    .Y(_03642_));
 sky130_fd_sc_hd__nand2_1 _09545_ (.A(_03540_),
    .B(_03543_),
    .Y(_03643_));
 sky130_fd_sc_hd__a31o_1 _09546_ (.A1(net398),
    .A2(net522),
    .A3(_03512_),
    .B1(_03511_),
    .X(_03644_));
 sky130_fd_sc_hd__nand4_1 _09547_ (.A(net390),
    .B(net374),
    .C(net530),
    .D(net525),
    .Y(_03645_));
 sky130_fd_sc_hd__a22o_1 _09548_ (.A1(net374),
    .A2(net530),
    .B1(net522),
    .B2(net390),
    .X(_03647_));
 sky130_fd_sc_hd__a22o_1 _09549_ (.A1(net365),
    .A2(net536),
    .B1(_03645_),
    .B2(_03647_),
    .X(_03648_));
 sky130_fd_sc_hd__nand4_1 _09550_ (.A(net365),
    .B(net537),
    .C(_03645_),
    .D(_03647_),
    .Y(_03649_));
 sky130_fd_sc_hd__nand3_1 _09551_ (.A(_03644_),
    .B(_03648_),
    .C(_03649_),
    .Y(_03650_));
 sky130_fd_sc_hd__a21o_1 _09552_ (.A1(_03648_),
    .A2(_03649_),
    .B1(_03644_),
    .X(_03651_));
 sky130_fd_sc_hd__nand3_1 _09553_ (.A(_03643_),
    .B(_03650_),
    .C(_03651_),
    .Y(_03652_));
 sky130_fd_sc_hd__a21o_1 _09554_ (.A1(_03650_),
    .A2(_03651_),
    .B1(_03643_),
    .X(_03653_));
 sky130_fd_sc_hd__a21bo_1 _09555_ (.A1(_03538_),
    .A2(_03545_),
    .B1_N(_03544_),
    .X(_03654_));
 sky130_fd_sc_hd__and3_1 _09556_ (.A(_03652_),
    .B(_03653_),
    .C(_03654_),
    .X(_03655_));
 sky130_fd_sc_hd__a21oi_1 _09557_ (.A1(_03652_),
    .A2(_03653_),
    .B1(_03654_),
    .Y(_03656_));
 sky130_fd_sc_hd__or3_1 _09558_ (.A(_03642_),
    .B(_03655_),
    .C(_03656_),
    .X(_03658_));
 sky130_fd_sc_hd__o21ai_1 _09559_ (.A1(_03655_),
    .A2(_03656_),
    .B1(_03642_),
    .Y(_03659_));
 sky130_fd_sc_hd__and3_1 _09560_ (.A(_03518_),
    .B(_03658_),
    .C(_03659_),
    .X(_03660_));
 sky130_fd_sc_hd__nand3_1 _09561_ (.A(_03518_),
    .B(_03658_),
    .C(_03659_),
    .Y(_03661_));
 sky130_fd_sc_hd__a21oi_1 _09562_ (.A1(_03658_),
    .A2(_03659_),
    .B1(_03518_),
    .Y(_03662_));
 sky130_fd_sc_hd__a211o_1 _09563_ (.A1(_03551_),
    .A2(_03553_),
    .B1(_03660_),
    .C1(_03662_),
    .X(_03663_));
 sky130_fd_sc_hd__o211ai_2 _09564_ (.A1(_03660_),
    .A2(_03662_),
    .B1(_03551_),
    .C1(_03553_),
    .Y(_03664_));
 sky130_fd_sc_hd__nand4_2 _09565_ (.A(_03623_),
    .B(_03626_),
    .C(_03663_),
    .D(_03664_),
    .Y(_03665_));
 sky130_fd_sc_hd__a22o_1 _09566_ (.A1(_03623_),
    .A2(_03626_),
    .B1(_03663_),
    .B2(_03664_),
    .X(_03666_));
 sky130_fd_sc_hd__a21oi_1 _09567_ (.A1(_03665_),
    .A2(_03666_),
    .B1(_03561_),
    .Y(_03667_));
 sky130_fd_sc_hd__and3_1 _09568_ (.A(_03561_),
    .B(_03665_),
    .C(_03666_),
    .X(_03669_));
 sky130_fd_sc_hd__inv_2 _09569_ (.A(_03669_),
    .Y(_03670_));
 sky130_fd_sc_hd__nand2_1 _09570_ (.A(_03598_),
    .B(_03600_),
    .Y(_03671_));
 sky130_fd_sc_hd__and4_1 _09571_ (.A(net167),
    .B(net159),
    .C(net275),
    .D(net266),
    .X(_03672_));
 sky130_fd_sc_hd__a22oi_1 _09572_ (.A1(net159),
    .A2(net275),
    .B1(net266),
    .B2(net167),
    .Y(_03673_));
 sky130_fd_sc_hd__o2bb2a_1 _09573_ (.A1_N(net175),
    .A2_N(net259),
    .B1(_03672_),
    .B2(_03673_),
    .X(_03674_));
 sky130_fd_sc_hd__and4bb_1 _09574_ (.A_N(_03672_),
    .B_N(_03673_),
    .C(net175),
    .D(net259),
    .X(_03675_));
 sky130_fd_sc_hd__nor2_1 _09575_ (.A(_03674_),
    .B(_03675_),
    .Y(_03676_));
 sky130_fd_sc_hd__nor2_1 _09576_ (.A(_03565_),
    .B(_03568_),
    .Y(_03677_));
 sky130_fd_sc_hd__and2b_1 _09577_ (.A_N(_03677_),
    .B(_03676_),
    .X(_03678_));
 sky130_fd_sc_hd__xnor2_1 _09578_ (.A(_03676_),
    .B(_03677_),
    .Y(_03680_));
 sky130_fd_sc_hd__nand2_1 _09579_ (.A(net220),
    .B(net249),
    .Y(_03681_));
 sky130_fd_sc_hd__inv_2 _09580_ (.A(_03681_),
    .Y(_03682_));
 sky130_fd_sc_hd__xnor2_1 _09581_ (.A(_03680_),
    .B(_03682_),
    .Y(_03683_));
 sky130_fd_sc_hd__a21oi_1 _09582_ (.A1(_03573_),
    .A2(_03574_),
    .B1(_03572_),
    .Y(_03684_));
 sky130_fd_sc_hd__or2_1 _09583_ (.A(_03683_),
    .B(_03684_),
    .X(_03685_));
 sky130_fd_sc_hd__xor2_1 _09584_ (.A(_03683_),
    .B(_03684_),
    .X(_03686_));
 sky130_fd_sc_hd__nand2_1 _09585_ (.A(net297),
    .B(net243),
    .Y(_03687_));
 sky130_fd_sc_hd__nand3_1 _09586_ (.A(net297),
    .B(net243),
    .C(_03686_),
    .Y(_03688_));
 sky130_fd_sc_hd__xnor2_1 _09587_ (.A(_03686_),
    .B(_03687_),
    .Y(_03689_));
 sky130_fd_sc_hd__a21o_1 _09588_ (.A1(_03525_),
    .A2(_03534_),
    .B1(_03533_),
    .X(_03691_));
 sky130_fd_sc_hd__nand2_1 _09589_ (.A(_03585_),
    .B(_03588_),
    .Y(_03692_));
 sky130_fd_sc_hd__a31o_1 _09590_ (.A1(net591),
    .A2(net312),
    .A3(_03522_),
    .B1(_03521_),
    .X(_03693_));
 sky130_fd_sc_hd__nand4_2 _09591_ (.A(net607),
    .B(net591),
    .C(net304),
    .D(net290),
    .Y(_03694_));
 sky130_fd_sc_hd__a22o_1 _09592_ (.A1(net591),
    .A2(net304),
    .B1(net290),
    .B2(net607),
    .X(_03695_));
 sky130_fd_sc_hd__a22o_1 _09593_ (.A1(net616),
    .A2(net283),
    .B1(_03694_),
    .B2(_03695_),
    .X(_03696_));
 sky130_fd_sc_hd__nand4_2 _09594_ (.A(net616),
    .B(net283),
    .C(_03694_),
    .D(_03695_),
    .Y(_03697_));
 sky130_fd_sc_hd__nand3_2 _09595_ (.A(_03693_),
    .B(_03696_),
    .C(_03697_),
    .Y(_03698_));
 sky130_fd_sc_hd__a21o_1 _09596_ (.A1(_03696_),
    .A2(_03697_),
    .B1(_03693_),
    .X(_03699_));
 sky130_fd_sc_hd__nand3_2 _09597_ (.A(_03692_),
    .B(_03698_),
    .C(_03699_),
    .Y(_03700_));
 sky130_fd_sc_hd__a21o_1 _09598_ (.A1(_03698_),
    .A2(_03699_),
    .B1(_03692_),
    .X(_03702_));
 sky130_fd_sc_hd__and3_1 _09599_ (.A(_03691_),
    .B(_03700_),
    .C(_03702_),
    .X(_03703_));
 sky130_fd_sc_hd__nand3_1 _09600_ (.A(_03691_),
    .B(_03700_),
    .C(_03702_),
    .Y(_03704_));
 sky130_fd_sc_hd__a21oi_1 _09601_ (.A1(_03700_),
    .A2(_03702_),
    .B1(_03691_),
    .Y(_03705_));
 sky130_fd_sc_hd__a211o_1 _09602_ (.A1(_03589_),
    .A2(_03591_),
    .B1(_03703_),
    .C1(_03705_),
    .X(_03706_));
 sky130_fd_sc_hd__o211ai_2 _09603_ (.A1(_03703_),
    .A2(_03705_),
    .B1(_03589_),
    .C1(_03591_),
    .Y(_03707_));
 sky130_fd_sc_hd__o211ai_2 _09604_ (.A1(_03594_),
    .A2(_03596_),
    .B1(_03706_),
    .C1(_03707_),
    .Y(_03708_));
 sky130_fd_sc_hd__a211o_1 _09605_ (.A1(_03706_),
    .A2(_03707_),
    .B1(_03594_),
    .C1(_03596_),
    .X(_03709_));
 sky130_fd_sc_hd__and3_1 _09606_ (.A(_03689_),
    .B(_03708_),
    .C(_03709_),
    .X(_03710_));
 sky130_fd_sc_hd__inv_2 _09607_ (.A(_03710_),
    .Y(_03711_));
 sky130_fd_sc_hd__a21oi_1 _09608_ (.A1(_03708_),
    .A2(_03709_),
    .B1(_03689_),
    .Y(_03713_));
 sky130_fd_sc_hd__a211o_1 _09609_ (.A1(_03556_),
    .A2(_03558_),
    .B1(_03710_),
    .C1(_03713_),
    .X(_03714_));
 sky130_fd_sc_hd__o211ai_1 _09610_ (.A1(_03710_),
    .A2(_03713_),
    .B1(_03556_),
    .C1(_03558_),
    .Y(_03715_));
 sky130_fd_sc_hd__and3_1 _09611_ (.A(_03671_),
    .B(_03714_),
    .C(_03715_),
    .X(_03716_));
 sky130_fd_sc_hd__inv_2 _09612_ (.A(_03716_),
    .Y(_03717_));
 sky130_fd_sc_hd__a21oi_1 _09613_ (.A1(_03714_),
    .A2(_03715_),
    .B1(_03671_),
    .Y(_03718_));
 sky130_fd_sc_hd__nor4_1 _09614_ (.A(_03667_),
    .B(_03669_),
    .C(_03716_),
    .D(_03718_),
    .Y(_03719_));
 sky130_fd_sc_hd__or4_1 _09615_ (.A(_03667_),
    .B(_03669_),
    .C(_03716_),
    .D(_03718_),
    .X(_03720_));
 sky130_fd_sc_hd__o22a_1 _09616_ (.A1(_03667_),
    .A2(_03669_),
    .B1(_03716_),
    .B2(_03718_),
    .X(_03721_));
 sky130_fd_sc_hd__a211oi_2 _09617_ (.A1(_03564_),
    .A2(_03608_),
    .B1(net134),
    .C1(_03721_),
    .Y(_03722_));
 sky130_fd_sc_hd__inv_2 _09618_ (.A(_03722_),
    .Y(_03724_));
 sky130_fd_sc_hd__o211a_1 _09619_ (.A1(_03719_),
    .A2(_03721_),
    .B1(_03564_),
    .C1(_03608_),
    .X(_03725_));
 sky130_fd_sc_hd__a211o_1 _09620_ (.A1(_03604_),
    .A2(_03606_),
    .B1(_03722_),
    .C1(_03725_),
    .X(_03726_));
 sky130_fd_sc_hd__o211ai_1 _09621_ (.A1(_03722_),
    .A2(_03725_),
    .B1(_03604_),
    .C1(_03606_),
    .Y(_03727_));
 sky130_fd_sc_hd__nand2_1 _09622_ (.A(_03726_),
    .B(_03727_),
    .Y(_03728_));
 sky130_fd_sc_hd__or2_1 _09623_ (.A(_03610_),
    .B(_03612_),
    .X(_03729_));
 sky130_fd_sc_hd__xnor2_1 _09624_ (.A(_03728_),
    .B(_03729_),
    .Y(_03730_));
 sky130_fd_sc_hd__o21ai_1 _09625_ (.A1(_03575_),
    .A2(_03576_),
    .B1(_03579_),
    .Y(_03731_));
 sky130_fd_sc_hd__xnor2_1 _09626_ (.A(_03730_),
    .B(_03731_),
    .Y(_03732_));
 sky130_fd_sc_hd__nor2_1 _09627_ (.A(_03615_),
    .B(_03617_),
    .Y(_03733_));
 sky130_fd_sc_hd__nor2_1 _09628_ (.A(_03732_),
    .B(_03733_),
    .Y(_03735_));
 sky130_fd_sc_hd__xor2_1 _09629_ (.A(_03732_),
    .B(_03733_),
    .X(_03736_));
 sky130_fd_sc_hd__o21ba_1 _09630_ (.A1(_03506_),
    .A2(_03620_),
    .B1_N(_03619_),
    .X(_03737_));
 sky130_fd_sc_hd__nand2_1 _09631_ (.A(_03508_),
    .B(_03621_),
    .Y(_03738_));
 sky130_fd_sc_hd__inv_2 _09632_ (.A(_03738_),
    .Y(_03739_));
 sky130_fd_sc_hd__a21oi_2 _09633_ (.A1(_03510_),
    .A2(_03739_),
    .B1(_03737_),
    .Y(_03740_));
 sky130_fd_sc_hd__and2b_1 _09634_ (.A_N(_03740_),
    .B(_03736_),
    .X(_03741_));
 sky130_fd_sc_hd__xnor2_1 _09635_ (.A(_03736_),
    .B(_03740_),
    .Y(net103));
 sky130_fd_sc_hd__and2_1 _09636_ (.A(net377),
    .B(net511),
    .X(_03742_));
 sky130_fd_sc_hd__nand2_1 _09637_ (.A(net377),
    .B(net511),
    .Y(_03743_));
 sky130_fd_sc_hd__and4_1 _09638_ (.A(net390),
    .B(net374),
    .C(net525),
    .D(net513),
    .X(_03745_));
 sky130_fd_sc_hd__a22oi_1 _09639_ (.A1(net374),
    .A2(net525),
    .B1(net513),
    .B2(net390),
    .Y(_03746_));
 sky130_fd_sc_hd__o2bb2a_1 _09640_ (.A1_N(net366),
    .A2_N(net531),
    .B1(_03745_),
    .B2(_03746_),
    .X(_03747_));
 sky130_fd_sc_hd__and4bb_1 _09641_ (.A_N(_03745_),
    .B_N(_03746_),
    .C(net366),
    .D(net531),
    .X(_03748_));
 sky130_fd_sc_hd__or3_1 _09642_ (.A(_03626_),
    .B(_03747_),
    .C(_03748_),
    .X(_03749_));
 sky130_fd_sc_hd__o21ai_1 _09643_ (.A1(_03747_),
    .A2(_03748_),
    .B1(_03626_),
    .Y(_03750_));
 sky130_fd_sc_hd__nand2_1 _09644_ (.A(_03645_),
    .B(_03649_),
    .Y(_03751_));
 sky130_fd_sc_hd__a21oi_1 _09645_ (.A1(_03749_),
    .A2(_03750_),
    .B1(_03751_),
    .Y(_03752_));
 sky130_fd_sc_hd__and3_1 _09646_ (.A(_03749_),
    .B(_03750_),
    .C(_03751_),
    .X(_03753_));
 sky130_fd_sc_hd__or2_1 _09647_ (.A(_03752_),
    .B(_03753_),
    .X(_03754_));
 sky130_fd_sc_hd__nand2_1 _09648_ (.A(_03650_),
    .B(_03652_),
    .Y(_03756_));
 sky130_fd_sc_hd__and2b_1 _09649_ (.A_N(_03754_),
    .B(_03756_),
    .X(_03757_));
 sky130_fd_sc_hd__xor2_1 _09650_ (.A(_03754_),
    .B(_03756_),
    .X(_03758_));
 sky130_fd_sc_hd__and4_1 _09651_ (.A(net328),
    .B(net320),
    .C(net571),
    .D(net564),
    .X(_03759_));
 sky130_fd_sc_hd__a22o_1 _09652_ (.A1(net320),
    .A2(net571),
    .B1(net564),
    .B2(net328),
    .X(_03760_));
 sky130_fd_sc_hd__and2b_1 _09653_ (.A_N(_03759_),
    .B(_03760_),
    .X(_03761_));
 sky130_fd_sc_hd__nand2_1 _09654_ (.A(net577),
    .B(net312),
    .Y(_03762_));
 sky130_fd_sc_hd__xnor2_1 _09655_ (.A(_03761_),
    .B(_03762_),
    .Y(_03763_));
 sky130_fd_sc_hd__nand4_1 _09656_ (.A(net358),
    .B(net350),
    .C(net550),
    .D(net537),
    .Y(_03764_));
 sky130_fd_sc_hd__a22o_1 _09657_ (.A1(net350),
    .A2(net550),
    .B1(net537),
    .B2(net358),
    .X(_03765_));
 sky130_fd_sc_hd__and2_1 _09658_ (.A(net335),
    .B(net557),
    .X(_03767_));
 sky130_fd_sc_hd__a21o_1 _09659_ (.A1(_03764_),
    .A2(_03765_),
    .B1(_03767_),
    .X(_03768_));
 sky130_fd_sc_hd__nand3_1 _09660_ (.A(_03764_),
    .B(_03765_),
    .C(_03767_),
    .Y(_03769_));
 sky130_fd_sc_hd__a21bo_1 _09661_ (.A1(_03633_),
    .A2(_03634_),
    .B1_N(_03632_),
    .X(_03770_));
 sky130_fd_sc_hd__and3_1 _09662_ (.A(_03768_),
    .B(_03769_),
    .C(_03770_),
    .X(_03771_));
 sky130_fd_sc_hd__a21o_1 _09663_ (.A1(_03768_),
    .A2(_03769_),
    .B1(_03770_),
    .X(_03772_));
 sky130_fd_sc_hd__and2b_1 _09664_ (.A_N(_03771_),
    .B(_03772_),
    .X(_03773_));
 sky130_fd_sc_hd__xnor2_1 _09665_ (.A(_03763_),
    .B(_03773_),
    .Y(_03774_));
 sky130_fd_sc_hd__nor2_1 _09666_ (.A(_03758_),
    .B(_03774_),
    .Y(_03775_));
 sky130_fd_sc_hd__xnor2_1 _09667_ (.A(_03758_),
    .B(_03774_),
    .Y(_03776_));
 sky130_fd_sc_hd__nand2b_1 _09668_ (.A_N(_03655_),
    .B(_03658_),
    .Y(_03778_));
 sky130_fd_sc_hd__and2b_1 _09669_ (.A_N(_03776_),
    .B(_03778_),
    .X(_03779_));
 sky130_fd_sc_hd__xnor2_1 _09670_ (.A(_03776_),
    .B(_03778_),
    .Y(_03780_));
 sky130_fd_sc_hd__nand2b_1 _09671_ (.A_N(_03625_),
    .B(_03780_),
    .Y(_03781_));
 sky130_fd_sc_hd__xnor2_1 _09672_ (.A(_03625_),
    .B(_03780_),
    .Y(_03782_));
 sky130_fd_sc_hd__and2b_1 _09673_ (.A_N(_03665_),
    .B(_03782_),
    .X(_03783_));
 sky130_fd_sc_hd__xnor2_1 _09674_ (.A(_03665_),
    .B(_03782_),
    .Y(_03784_));
 sky130_fd_sc_hd__and4_1 _09675_ (.A(net159),
    .B(net615),
    .C(net275),
    .D(net266),
    .X(_03785_));
 sky130_fd_sc_hd__a22oi_1 _09676_ (.A1(net615),
    .A2(net275),
    .B1(net266),
    .B2(net159),
    .Y(_03786_));
 sky130_fd_sc_hd__o2bb2a_1 _09677_ (.A1_N(net167),
    .A2_N(net259),
    .B1(_03785_),
    .B2(_03786_),
    .X(_03787_));
 sky130_fd_sc_hd__and4bb_1 _09678_ (.A_N(_03785_),
    .B_N(_03786_),
    .C(net167),
    .D(net259),
    .X(_03789_));
 sky130_fd_sc_hd__nor2_1 _09679_ (.A(_03787_),
    .B(_03789_),
    .Y(_03790_));
 sky130_fd_sc_hd__nor2_1 _09680_ (.A(_03672_),
    .B(_03675_),
    .Y(_03791_));
 sky130_fd_sc_hd__and2b_1 _09681_ (.A_N(_03791_),
    .B(_03790_),
    .X(_03792_));
 sky130_fd_sc_hd__xnor2_1 _09682_ (.A(_03790_),
    .B(_03791_),
    .Y(_03793_));
 sky130_fd_sc_hd__and2_1 _09683_ (.A(net175),
    .B(net249),
    .X(_03794_));
 sky130_fd_sc_hd__xnor2_1 _09684_ (.A(_03793_),
    .B(_03794_),
    .Y(_03795_));
 sky130_fd_sc_hd__a21oi_1 _09685_ (.A1(_03680_),
    .A2(_03682_),
    .B1(_03678_),
    .Y(_03796_));
 sky130_fd_sc_hd__xnor2_1 _09686_ (.A(_03795_),
    .B(_03796_),
    .Y(_03797_));
 sky130_fd_sc_hd__nand2_1 _09687_ (.A(net220),
    .B(net243),
    .Y(_03798_));
 sky130_fd_sc_hd__or2_1 _09688_ (.A(_03797_),
    .B(_03798_),
    .X(_03800_));
 sky130_fd_sc_hd__xor2_1 _09689_ (.A(_03797_),
    .B(_03798_),
    .X(_03801_));
 sky130_fd_sc_hd__a21o_1 _09690_ (.A1(_03631_),
    .A2(_03640_),
    .B1(_03639_),
    .X(_03802_));
 sky130_fd_sc_hd__nand2_1 _09691_ (.A(_03694_),
    .B(_03697_),
    .Y(_03803_));
 sky130_fd_sc_hd__a31o_1 _09692_ (.A1(net584),
    .A2(net313),
    .A3(_03628_),
    .B1(_03627_),
    .X(_03804_));
 sky130_fd_sc_hd__nand4_2 _09693_ (.A(net591),
    .B(net584),
    .C(net304),
    .D(net291),
    .Y(_03805_));
 sky130_fd_sc_hd__a22o_1 _09694_ (.A1(net584),
    .A2(net305),
    .B1(net291),
    .B2(net591),
    .X(_03806_));
 sky130_fd_sc_hd__a22o_1 _09695_ (.A1(net608),
    .A2(net284),
    .B1(_03805_),
    .B2(_03806_),
    .X(_03807_));
 sky130_fd_sc_hd__nand4_2 _09696_ (.A(net608),
    .B(net284),
    .C(_03805_),
    .D(_03806_),
    .Y(_03808_));
 sky130_fd_sc_hd__nand3_2 _09697_ (.A(_03804_),
    .B(_03807_),
    .C(_03808_),
    .Y(_03809_));
 sky130_fd_sc_hd__a21o_1 _09698_ (.A1(_03807_),
    .A2(_03808_),
    .B1(_03804_),
    .X(_03811_));
 sky130_fd_sc_hd__nand3_2 _09699_ (.A(_03803_),
    .B(_03809_),
    .C(_03811_),
    .Y(_03812_));
 sky130_fd_sc_hd__a21o_1 _09700_ (.A1(_03809_),
    .A2(_03811_),
    .B1(_03803_),
    .X(_03813_));
 sky130_fd_sc_hd__and3_2 _09701_ (.A(_03802_),
    .B(_03812_),
    .C(_03813_),
    .X(_03814_));
 sky130_fd_sc_hd__a21oi_2 _09702_ (.A1(_03812_),
    .A2(_03813_),
    .B1(_03802_),
    .Y(_03815_));
 sky130_fd_sc_hd__a211oi_4 _09703_ (.A1(_03698_),
    .A2(_03700_),
    .B1(_03814_),
    .C1(_03815_),
    .Y(_03816_));
 sky130_fd_sc_hd__o211a_1 _09704_ (.A1(_03814_),
    .A2(_03815_),
    .B1(_03698_),
    .C1(_03700_),
    .X(_03817_));
 sky130_fd_sc_hd__a211o_1 _09705_ (.A1(_03704_),
    .A2(_03706_),
    .B1(_03816_),
    .C1(_03817_),
    .X(_03818_));
 sky130_fd_sc_hd__inv_2 _09706_ (.A(_03818_),
    .Y(_03819_));
 sky130_fd_sc_hd__o211ai_1 _09707_ (.A1(_03816_),
    .A2(_03817_),
    .B1(_03704_),
    .C1(_03706_),
    .Y(_03820_));
 sky130_fd_sc_hd__and3_2 _09708_ (.A(_03801_),
    .B(_03818_),
    .C(_03820_),
    .X(_03822_));
 sky130_fd_sc_hd__a21oi_1 _09709_ (.A1(_03818_),
    .A2(_03820_),
    .B1(_03801_),
    .Y(_03823_));
 sky130_fd_sc_hd__a211oi_1 _09710_ (.A1(_03661_),
    .A2(_03663_),
    .B1(_03822_),
    .C1(_03823_),
    .Y(_03824_));
 sky130_fd_sc_hd__a211o_1 _09711_ (.A1(_03661_),
    .A2(_03663_),
    .B1(_03822_),
    .C1(_03823_),
    .X(_03825_));
 sky130_fd_sc_hd__o211a_1 _09712_ (.A1(_03822_),
    .A2(_03823_),
    .B1(_03661_),
    .C1(_03663_),
    .X(_03826_));
 sky130_fd_sc_hd__a211o_1 _09713_ (.A1(_03708_),
    .A2(_03711_),
    .B1(_03824_),
    .C1(_03826_),
    .X(_03827_));
 sky130_fd_sc_hd__o211ai_1 _09714_ (.A1(_03824_),
    .A2(_03826_),
    .B1(_03708_),
    .C1(_03711_),
    .Y(_03828_));
 sky130_fd_sc_hd__and3_1 _09715_ (.A(_03784_),
    .B(_03827_),
    .C(_03828_),
    .X(_03829_));
 sky130_fd_sc_hd__a21oi_1 _09716_ (.A1(_03827_),
    .A2(_03828_),
    .B1(_03784_),
    .Y(_03830_));
 sky130_fd_sc_hd__a211oi_2 _09717_ (.A1(_03670_),
    .A2(_03720_),
    .B1(_03829_),
    .C1(_03830_),
    .Y(_03831_));
 sky130_fd_sc_hd__o211a_1 _09718_ (.A1(_03829_),
    .A2(_03830_),
    .B1(_03670_),
    .C1(_03720_),
    .X(_03833_));
 sky130_fd_sc_hd__a211oi_2 _09719_ (.A1(_03714_),
    .A2(_03717_),
    .B1(_03831_),
    .C1(_03833_),
    .Y(_03834_));
 sky130_fd_sc_hd__o211a_1 _09720_ (.A1(_03831_),
    .A2(_03833_),
    .B1(_03714_),
    .C1(_03717_),
    .X(_03835_));
 sky130_fd_sc_hd__a211oi_1 _09721_ (.A1(_03724_),
    .A2(_03726_),
    .B1(_03834_),
    .C1(_03835_),
    .Y(_03836_));
 sky130_fd_sc_hd__o211a_1 _09722_ (.A1(_03834_),
    .A2(_03835_),
    .B1(_03724_),
    .C1(_03726_),
    .X(_03837_));
 sky130_fd_sc_hd__a211o_1 _09723_ (.A1(_03685_),
    .A2(_03688_),
    .B1(_03836_),
    .C1(_03837_),
    .X(_03838_));
 sky130_fd_sc_hd__o211ai_1 _09724_ (.A1(_03836_),
    .A2(_03837_),
    .B1(_03685_),
    .C1(_03688_),
    .Y(_03839_));
 sky130_fd_sc_hd__nand2_1 _09725_ (.A(_03838_),
    .B(_03839_),
    .Y(_03840_));
 sky130_fd_sc_hd__a32o_1 _09726_ (.A1(_03726_),
    .A2(_03727_),
    .A3(_03729_),
    .B1(_03730_),
    .B2(_03731_),
    .X(_03841_));
 sky130_fd_sc_hd__nand2b_1 _09727_ (.A_N(_03841_),
    .B(_03840_),
    .Y(_03842_));
 sky130_fd_sc_hd__and3_1 _09728_ (.A(_03838_),
    .B(_03839_),
    .C(_03841_),
    .X(_03844_));
 sky130_fd_sc_hd__xnor2_1 _09729_ (.A(_03840_),
    .B(_03841_),
    .Y(_03845_));
 sky130_fd_sc_hd__nor2_1 _09730_ (.A(_03735_),
    .B(_03741_),
    .Y(_03846_));
 sky130_fd_sc_hd__xnor2_1 _09731_ (.A(_03845_),
    .B(_03846_),
    .Y(net104));
 sky130_fd_sc_hd__and3_1 _09732_ (.A(net393),
    .B(net504),
    .C(_03742_),
    .X(_03847_));
 sky130_fd_sc_hd__a21o_1 _09733_ (.A1(net393),
    .A2(net504),
    .B1(_03742_),
    .X(_03848_));
 sky130_fd_sc_hd__and2b_1 _09734_ (.A_N(_03847_),
    .B(_03848_),
    .X(_03849_));
 sky130_fd_sc_hd__nand2_1 _09735_ (.A(net367),
    .B(net525),
    .Y(_03850_));
 sky130_fd_sc_hd__xnor2_1 _09736_ (.A(_03849_),
    .B(_03850_),
    .Y(_03851_));
 sky130_fd_sc_hd__nor2_1 _09737_ (.A(_03745_),
    .B(_03748_),
    .Y(_03852_));
 sky130_fd_sc_hd__and2b_1 _09738_ (.A_N(_03852_),
    .B(_03851_),
    .X(_03854_));
 sky130_fd_sc_hd__xnor2_1 _09739_ (.A(_03851_),
    .B(_03852_),
    .Y(_03855_));
 sky130_fd_sc_hd__a21boi_1 _09740_ (.A1(_03750_),
    .A2(_03751_),
    .B1_N(_03749_),
    .Y(_03856_));
 sky130_fd_sc_hd__nand2b_1 _09741_ (.A_N(_03856_),
    .B(_03855_),
    .Y(_03857_));
 sky130_fd_sc_hd__xnor2_1 _09742_ (.A(_03855_),
    .B(_03856_),
    .Y(_03858_));
 sky130_fd_sc_hd__and4_1 _09743_ (.A(net328),
    .B(net320),
    .C(net567),
    .D(net560),
    .X(_03859_));
 sky130_fd_sc_hd__a22o_1 _09744_ (.A1(net322),
    .A2(net567),
    .B1(net560),
    .B2(net329),
    .X(_03860_));
 sky130_fd_sc_hd__and2b_1 _09745_ (.A_N(_03859_),
    .B(_03860_),
    .X(_03861_));
 sky130_fd_sc_hd__nand2_1 _09746_ (.A(net574),
    .B(net313),
    .Y(_03862_));
 sky130_fd_sc_hd__xnor2_1 _09747_ (.A(_03861_),
    .B(_03862_),
    .Y(_03863_));
 sky130_fd_sc_hd__nand4_1 _09748_ (.A(net358),
    .B(net350),
    .C(net539),
    .D(net531),
    .Y(_03865_));
 sky130_fd_sc_hd__a22o_1 _09749_ (.A1(net351),
    .A2(net539),
    .B1(net533),
    .B2(net359),
    .X(_03866_));
 sky130_fd_sc_hd__a22o_1 _09750_ (.A1(net335),
    .A2(net555),
    .B1(_03865_),
    .B2(_03866_),
    .X(_03867_));
 sky130_fd_sc_hd__nand4_1 _09751_ (.A(net336),
    .B(net555),
    .C(_03865_),
    .D(_03866_),
    .Y(_03868_));
 sky130_fd_sc_hd__a21bo_1 _09752_ (.A1(_03765_),
    .A2(_03767_),
    .B1_N(_03764_),
    .X(_03869_));
 sky130_fd_sc_hd__and3_1 _09753_ (.A(_03867_),
    .B(_03868_),
    .C(_03869_),
    .X(_03870_));
 sky130_fd_sc_hd__a21o_1 _09754_ (.A1(_03867_),
    .A2(_03868_),
    .B1(_03869_),
    .X(_03871_));
 sky130_fd_sc_hd__and2b_1 _09755_ (.A_N(_03870_),
    .B(_03871_),
    .X(_03872_));
 sky130_fd_sc_hd__xnor2_1 _09756_ (.A(_03863_),
    .B(_03872_),
    .Y(_03873_));
 sky130_fd_sc_hd__inv_2 _09757_ (.A(_03873_),
    .Y(_03874_));
 sky130_fd_sc_hd__nand2_1 _09758_ (.A(_03858_),
    .B(_03874_),
    .Y(_03876_));
 sky130_fd_sc_hd__xnor2_1 _09759_ (.A(_03858_),
    .B(_03874_),
    .Y(_03877_));
 sky130_fd_sc_hd__o21ba_1 _09760_ (.A1(_03757_),
    .A2(_03775_),
    .B1_N(_03877_),
    .X(_03878_));
 sky130_fd_sc_hd__or3b_1 _09761_ (.A(_03757_),
    .B(_03775_),
    .C_N(_03877_),
    .X(_03879_));
 sky130_fd_sc_hd__nand2b_1 _09762_ (.A_N(_03878_),
    .B(_03879_),
    .Y(_03880_));
 sky130_fd_sc_hd__nand2_1 _09763_ (.A(_03781_),
    .B(_03880_),
    .Y(_03881_));
 sky130_fd_sc_hd__or2_1 _09764_ (.A(_03781_),
    .B(_03880_),
    .X(_03882_));
 sky130_fd_sc_hd__inv_2 _09765_ (.A(_03882_),
    .Y(_03883_));
 sky130_fd_sc_hd__and4_1 _09766_ (.A(net615),
    .B(net607),
    .C(net275),
    .D(net266),
    .X(_03884_));
 sky130_fd_sc_hd__a22oi_1 _09767_ (.A1(net607),
    .A2(net275),
    .B1(net266),
    .B2(net615),
    .Y(_03885_));
 sky130_fd_sc_hd__o2bb2a_1 _09768_ (.A1_N(net160),
    .A2_N(net259),
    .B1(_03884_),
    .B2(_03885_),
    .X(_03887_));
 sky130_fd_sc_hd__and4bb_1 _09769_ (.A_N(_03884_),
    .B_N(_03885_),
    .C(net160),
    .D(net259),
    .X(_03888_));
 sky130_fd_sc_hd__nor2_1 _09770_ (.A(_03887_),
    .B(_03888_),
    .Y(_03889_));
 sky130_fd_sc_hd__nor2_1 _09771_ (.A(_03785_),
    .B(_03789_),
    .Y(_03890_));
 sky130_fd_sc_hd__and2b_1 _09772_ (.A_N(_03890_),
    .B(_03889_),
    .X(_03891_));
 sky130_fd_sc_hd__xnor2_1 _09773_ (.A(_03889_),
    .B(_03890_),
    .Y(_03892_));
 sky130_fd_sc_hd__and2_1 _09774_ (.A(net168),
    .B(net249),
    .X(_03893_));
 sky130_fd_sc_hd__xnor2_1 _09775_ (.A(_03892_),
    .B(_03893_),
    .Y(_03894_));
 sky130_fd_sc_hd__a21oi_1 _09776_ (.A1(_03793_),
    .A2(_03794_),
    .B1(_03792_),
    .Y(_03895_));
 sky130_fd_sc_hd__or2_1 _09777_ (.A(_03894_),
    .B(_03895_),
    .X(_03896_));
 sky130_fd_sc_hd__xnor2_1 _09778_ (.A(_03894_),
    .B(_03895_),
    .Y(_03898_));
 sky130_fd_sc_hd__nand2_1 _09779_ (.A(net176),
    .B(net243),
    .Y(_03899_));
 sky130_fd_sc_hd__or2_1 _09780_ (.A(_03898_),
    .B(_03899_),
    .X(_03900_));
 sky130_fd_sc_hd__xor2_1 _09781_ (.A(_03898_),
    .B(_03899_),
    .X(_03901_));
 sky130_fd_sc_hd__a21o_1 _09782_ (.A1(_03763_),
    .A2(_03772_),
    .B1(_03771_),
    .X(_03902_));
 sky130_fd_sc_hd__nand2_1 _09783_ (.A(_03805_),
    .B(_03808_),
    .Y(_03903_));
 sky130_fd_sc_hd__a31o_1 _09784_ (.A1(net577),
    .A2(net313),
    .A3(_03760_),
    .B1(_03759_),
    .X(_03904_));
 sky130_fd_sc_hd__nand4_2 _09785_ (.A(net585),
    .B(net578),
    .C(net306),
    .D(net291),
    .Y(_03905_));
 sky130_fd_sc_hd__a22o_1 _09786_ (.A1(net578),
    .A2(net306),
    .B1(net291),
    .B2(net585),
    .X(_03906_));
 sky130_fd_sc_hd__a22o_1 _09787_ (.A1(net592),
    .A2(net284),
    .B1(_03905_),
    .B2(_03906_),
    .X(_03907_));
 sky130_fd_sc_hd__nand4_2 _09788_ (.A(net592),
    .B(net284),
    .C(_03905_),
    .D(_03906_),
    .Y(_03909_));
 sky130_fd_sc_hd__nand3_2 _09789_ (.A(_03904_),
    .B(_03907_),
    .C(_03909_),
    .Y(_03910_));
 sky130_fd_sc_hd__a21o_1 _09790_ (.A1(_03907_),
    .A2(_03909_),
    .B1(_03904_),
    .X(_03911_));
 sky130_fd_sc_hd__nand3_2 _09791_ (.A(_03903_),
    .B(_03910_),
    .C(_03911_),
    .Y(_03912_));
 sky130_fd_sc_hd__a21o_1 _09792_ (.A1(_03910_),
    .A2(_03911_),
    .B1(_03903_),
    .X(_03913_));
 sky130_fd_sc_hd__and3_1 _09793_ (.A(_03902_),
    .B(_03912_),
    .C(_03913_),
    .X(_03914_));
 sky130_fd_sc_hd__nand3_1 _09794_ (.A(_03902_),
    .B(_03912_),
    .C(_03913_),
    .Y(_03915_));
 sky130_fd_sc_hd__a21oi_1 _09795_ (.A1(_03912_),
    .A2(_03913_),
    .B1(_03902_),
    .Y(_03916_));
 sky130_fd_sc_hd__a211o_2 _09796_ (.A1(_03809_),
    .A2(_03812_),
    .B1(_03914_),
    .C1(_03916_),
    .X(_03917_));
 sky130_fd_sc_hd__o211ai_2 _09797_ (.A1(_03914_),
    .A2(_03916_),
    .B1(_03809_),
    .C1(_03812_),
    .Y(_03918_));
 sky130_fd_sc_hd__o211ai_4 _09798_ (.A1(_03814_),
    .A2(_03816_),
    .B1(_03917_),
    .C1(_03918_),
    .Y(_03920_));
 sky130_fd_sc_hd__a211o_1 _09799_ (.A1(_03917_),
    .A2(_03918_),
    .B1(_03814_),
    .C1(_03816_),
    .X(_03921_));
 sky130_fd_sc_hd__nand3_2 _09800_ (.A(_03901_),
    .B(_03920_),
    .C(_03921_),
    .Y(_03922_));
 sky130_fd_sc_hd__a21o_1 _09801_ (.A1(_03920_),
    .A2(_03921_),
    .B1(_03901_),
    .X(_03923_));
 sky130_fd_sc_hd__nand3_2 _09802_ (.A(_03779_),
    .B(_03922_),
    .C(_03923_),
    .Y(_03924_));
 sky130_fd_sc_hd__a21o_1 _09803_ (.A1(_03922_),
    .A2(_03923_),
    .B1(_03779_),
    .X(_03925_));
 sky130_fd_sc_hd__o211ai_4 _09804_ (.A1(_03819_),
    .A2(_03822_),
    .B1(_03924_),
    .C1(_03925_),
    .Y(_03926_));
 sky130_fd_sc_hd__a211o_1 _09805_ (.A1(_03924_),
    .A2(_03925_),
    .B1(_03819_),
    .C1(_03822_),
    .X(_03927_));
 sky130_fd_sc_hd__and4_1 _09806_ (.A(_03881_),
    .B(_03882_),
    .C(_03926_),
    .D(_03927_),
    .X(_03928_));
 sky130_fd_sc_hd__nand4_1 _09807_ (.A(_03881_),
    .B(_03882_),
    .C(_03926_),
    .D(_03927_),
    .Y(_03929_));
 sky130_fd_sc_hd__a22o_1 _09808_ (.A1(_03881_),
    .A2(_03882_),
    .B1(_03926_),
    .B2(_03927_),
    .X(_03931_));
 sky130_fd_sc_hd__o211a_1 _09809_ (.A1(_03783_),
    .A2(_03829_),
    .B1(_03929_),
    .C1(_03931_),
    .X(_03932_));
 sky130_fd_sc_hd__inv_2 _09810_ (.A(_03932_),
    .Y(_03933_));
 sky130_fd_sc_hd__a211oi_1 _09811_ (.A1(_03929_),
    .A2(_03931_),
    .B1(_03783_),
    .C1(_03829_),
    .Y(_03934_));
 sky130_fd_sc_hd__a211o_1 _09812_ (.A1(_03825_),
    .A2(_03827_),
    .B1(_03932_),
    .C1(_03934_),
    .X(_03935_));
 sky130_fd_sc_hd__o211ai_2 _09813_ (.A1(_03932_),
    .A2(_03934_),
    .B1(_03825_),
    .C1(_03827_),
    .Y(_03936_));
 sky130_fd_sc_hd__o211a_1 _09814_ (.A1(_03831_),
    .A2(_03834_),
    .B1(_03935_),
    .C1(_03936_),
    .X(_03937_));
 sky130_fd_sc_hd__inv_2 _09815_ (.A(_03937_),
    .Y(_03938_));
 sky130_fd_sc_hd__a211oi_1 _09816_ (.A1(_03935_),
    .A2(_03936_),
    .B1(_03831_),
    .C1(_03834_),
    .Y(_03939_));
 sky130_fd_sc_hd__o21a_1 _09817_ (.A1(_03795_),
    .A2(_03796_),
    .B1(_03800_),
    .X(_03940_));
 sky130_fd_sc_hd__or3_1 _09818_ (.A(_03937_),
    .B(_03939_),
    .C(_03940_),
    .X(_03942_));
 sky130_fd_sc_hd__o21ai_1 _09819_ (.A1(_03937_),
    .A2(_03939_),
    .B1(_03940_),
    .Y(_03943_));
 sky130_fd_sc_hd__nand2_1 _09820_ (.A(_03942_),
    .B(_03943_),
    .Y(_03944_));
 sky130_fd_sc_hd__and2b_1 _09821_ (.A_N(_03836_),
    .B(_03838_),
    .X(_03945_));
 sky130_fd_sc_hd__nor2_1 _09822_ (.A(_03944_),
    .B(_03945_),
    .Y(_03946_));
 sky130_fd_sc_hd__xor2_1 _09823_ (.A(_03944_),
    .B(_03945_),
    .X(_03947_));
 sky130_fd_sc_hd__a21oi_1 _09824_ (.A1(_03735_),
    .A2(_03842_),
    .B1(_03844_),
    .Y(_03948_));
 sky130_fd_sc_hd__nand2_1 _09825_ (.A(_03736_),
    .B(_03845_),
    .Y(_03949_));
 sky130_fd_sc_hd__o21ai_1 _09826_ (.A1(_03740_),
    .A2(_03949_),
    .B1(_03948_),
    .Y(_03950_));
 sky130_fd_sc_hd__xor2_1 _09827_ (.A(_03947_),
    .B(_03950_),
    .X(net105));
 sky130_fd_sc_hd__a22o_1 _09828_ (.A1(net367),
    .A2(net511),
    .B1(net504),
    .B2(net377),
    .X(_03952_));
 sky130_fd_sc_hd__nand2_1 _09829_ (.A(net367),
    .B(net504),
    .Y(_03953_));
 sky130_fd_sc_hd__o21a_1 _09830_ (.A1(_03743_),
    .A2(_03953_),
    .B1(_03952_),
    .X(_03954_));
 sky130_fd_sc_hd__a31o_1 _09831_ (.A1(net367),
    .A2(net527),
    .A3(_03848_),
    .B1(_03847_),
    .X(_03955_));
 sky130_fd_sc_hd__nand2_1 _09832_ (.A(_03954_),
    .B(_03955_),
    .Y(_03956_));
 sky130_fd_sc_hd__or2_1 _09833_ (.A(_03954_),
    .B(_03955_),
    .X(_03957_));
 sky130_fd_sc_hd__and2_1 _09834_ (.A(_03956_),
    .B(_03957_),
    .X(_03958_));
 sky130_fd_sc_hd__nand2_1 _09835_ (.A(_03854_),
    .B(_03958_),
    .Y(_03959_));
 sky130_fd_sc_hd__xnor2_1 _09836_ (.A(_03854_),
    .B(_03958_),
    .Y(_03960_));
 sky130_fd_sc_hd__and4_1 _09837_ (.A(net329),
    .B(net322),
    .C(net561),
    .D(net555),
    .X(_03961_));
 sky130_fd_sc_hd__a22o_1 _09838_ (.A1(net322),
    .A2(net561),
    .B1(net555),
    .B2(net329),
    .X(_03963_));
 sky130_fd_sc_hd__and2b_1 _09839_ (.A_N(_03961_),
    .B(_03963_),
    .X(_03964_));
 sky130_fd_sc_hd__nand2_1 _09840_ (.A(net314),
    .B(net569),
    .Y(_03965_));
 sky130_fd_sc_hd__xnor2_1 _09841_ (.A(_03964_),
    .B(_03965_),
    .Y(_03966_));
 sky130_fd_sc_hd__nand4_1 _09842_ (.A(net359),
    .B(net351),
    .C(net534),
    .D(net524),
    .Y(_03967_));
 sky130_fd_sc_hd__a22o_1 _09843_ (.A1(net351),
    .A2(net534),
    .B1(net524),
    .B2(net359),
    .X(_03968_));
 sky130_fd_sc_hd__a22o_1 _09844_ (.A1(net336),
    .A2(net540),
    .B1(_03967_),
    .B2(_03968_),
    .X(_03969_));
 sky130_fd_sc_hd__nand4_1 _09845_ (.A(net336),
    .B(net540),
    .C(_03967_),
    .D(_03968_),
    .Y(_03970_));
 sky130_fd_sc_hd__nand2_1 _09846_ (.A(_03865_),
    .B(_03868_),
    .Y(_03971_));
 sky130_fd_sc_hd__and3_1 _09847_ (.A(_03969_),
    .B(_03970_),
    .C(_03971_),
    .X(_03972_));
 sky130_fd_sc_hd__a21o_1 _09848_ (.A1(_03969_),
    .A2(_03970_),
    .B1(_03971_),
    .X(_03974_));
 sky130_fd_sc_hd__and2b_1 _09849_ (.A_N(_03972_),
    .B(_03974_),
    .X(_03975_));
 sky130_fd_sc_hd__xnor2_1 _09850_ (.A(_03966_),
    .B(_03975_),
    .Y(_03976_));
 sky130_fd_sc_hd__nand2_1 _09851_ (.A(_03960_),
    .B(_03976_),
    .Y(_03977_));
 sky130_fd_sc_hd__or2_1 _09852_ (.A(_03960_),
    .B(_03976_),
    .X(_03978_));
 sky130_fd_sc_hd__nand2_1 _09853_ (.A(_03977_),
    .B(_03978_),
    .Y(_03979_));
 sky130_fd_sc_hd__a21oi_1 _09854_ (.A1(_03857_),
    .A2(_03876_),
    .B1(_03979_),
    .Y(_03980_));
 sky130_fd_sc_hd__and3_1 _09855_ (.A(_03857_),
    .B(_03876_),
    .C(_03979_),
    .X(_03981_));
 sky130_fd_sc_hd__or2_1 _09856_ (.A(_03980_),
    .B(_03981_),
    .X(_03982_));
 sky130_fd_sc_hd__and4_1 _09857_ (.A(net609),
    .B(net592),
    .C(net279),
    .D(net271),
    .X(_03983_));
 sky130_fd_sc_hd__a22oi_1 _09858_ (.A1(net592),
    .A2(net279),
    .B1(net271),
    .B2(net609),
    .Y(_03984_));
 sky130_fd_sc_hd__o2bb2a_1 _09859_ (.A1_N(net617),
    .A2_N(net261),
    .B1(_03983_),
    .B2(_03984_),
    .X(_03985_));
 sky130_fd_sc_hd__and4bb_1 _09860_ (.A_N(_03983_),
    .B_N(_03984_),
    .C(net617),
    .D(net261),
    .X(_03986_));
 sky130_fd_sc_hd__nor2_1 _09861_ (.A(_03985_),
    .B(_03986_),
    .Y(_03987_));
 sky130_fd_sc_hd__nor2_1 _09862_ (.A(_03884_),
    .B(_03888_),
    .Y(_03988_));
 sky130_fd_sc_hd__and2b_1 _09863_ (.A_N(_03988_),
    .B(_03987_),
    .X(_03989_));
 sky130_fd_sc_hd__xnor2_1 _09864_ (.A(_03987_),
    .B(_03988_),
    .Y(_03990_));
 sky130_fd_sc_hd__and2_1 _09865_ (.A(net166),
    .B(net251),
    .X(_03991_));
 sky130_fd_sc_hd__xnor2_1 _09866_ (.A(_03990_),
    .B(_03991_),
    .Y(_03992_));
 sky130_fd_sc_hd__a21oi_2 _09867_ (.A1(_03892_),
    .A2(_03893_),
    .B1(_03891_),
    .Y(_03993_));
 sky130_fd_sc_hd__xnor2_1 _09868_ (.A(_03992_),
    .B(_03993_),
    .Y(_03995_));
 sky130_fd_sc_hd__nand2_1 _09869_ (.A(net174),
    .B(net244),
    .Y(_03996_));
 sky130_fd_sc_hd__or2_1 _09870_ (.A(_03995_),
    .B(_03996_),
    .X(_03997_));
 sky130_fd_sc_hd__xor2_1 _09871_ (.A(_03995_),
    .B(_03996_),
    .X(_03998_));
 sky130_fd_sc_hd__a21o_1 _09872_ (.A1(_03863_),
    .A2(_03871_),
    .B1(_03870_),
    .X(_03999_));
 sky130_fd_sc_hd__nand2_1 _09873_ (.A(_03905_),
    .B(_03909_),
    .Y(_04000_));
 sky130_fd_sc_hd__a31o_1 _09874_ (.A1(net574),
    .A2(net315),
    .A3(_03860_),
    .B1(_03859_),
    .X(_04001_));
 sky130_fd_sc_hd__nand4_2 _09875_ (.A(net582),
    .B(net576),
    .C(net307),
    .D(net292),
    .Y(_04002_));
 sky130_fd_sc_hd__a22o_1 _09876_ (.A1(net576),
    .A2(net307),
    .B1(net292),
    .B2(net578),
    .X(_04003_));
 sky130_fd_sc_hd__a22o_1 _09877_ (.A1(net586),
    .A2(net285),
    .B1(_04002_),
    .B2(_04003_),
    .X(_04004_));
 sky130_fd_sc_hd__nand4_2 _09878_ (.A(net586),
    .B(net285),
    .C(_04002_),
    .D(_04003_),
    .Y(_04006_));
 sky130_fd_sc_hd__nand3_2 _09879_ (.A(_04001_),
    .B(_04004_),
    .C(_04006_),
    .Y(_04007_));
 sky130_fd_sc_hd__a21o_1 _09880_ (.A1(_04004_),
    .A2(_04006_),
    .B1(_04001_),
    .X(_04008_));
 sky130_fd_sc_hd__nand3_2 _09881_ (.A(_04000_),
    .B(_04007_),
    .C(_04008_),
    .Y(_04009_));
 sky130_fd_sc_hd__a21o_1 _09882_ (.A1(_04007_),
    .A2(_04008_),
    .B1(_04000_),
    .X(_04010_));
 sky130_fd_sc_hd__and3_1 _09883_ (.A(_03999_),
    .B(_04009_),
    .C(_04010_),
    .X(_04011_));
 sky130_fd_sc_hd__a21oi_1 _09884_ (.A1(_04009_),
    .A2(_04010_),
    .B1(_03999_),
    .Y(_04012_));
 sky130_fd_sc_hd__a211oi_2 _09885_ (.A1(_03910_),
    .A2(_03912_),
    .B1(_04011_),
    .C1(_04012_),
    .Y(_04013_));
 sky130_fd_sc_hd__o211a_1 _09886_ (.A1(_04011_),
    .A2(_04012_),
    .B1(_03910_),
    .C1(_03912_),
    .X(_04014_));
 sky130_fd_sc_hd__a211o_1 _09887_ (.A1(_03915_),
    .A2(_03917_),
    .B1(_04013_),
    .C1(_04014_),
    .X(_04015_));
 sky130_fd_sc_hd__o211ai_1 _09888_ (.A1(_04013_),
    .A2(_04014_),
    .B1(_03915_),
    .C1(_03917_),
    .Y(_04017_));
 sky130_fd_sc_hd__nand3_1 _09889_ (.A(_03998_),
    .B(_04015_),
    .C(_04017_),
    .Y(_04018_));
 sky130_fd_sc_hd__a21o_1 _09890_ (.A1(_04015_),
    .A2(_04017_),
    .B1(_03998_),
    .X(_04019_));
 sky130_fd_sc_hd__and3_1 _09891_ (.A(_03878_),
    .B(_04018_),
    .C(_04019_),
    .X(_04020_));
 sky130_fd_sc_hd__a21oi_1 _09892_ (.A1(_04018_),
    .A2(_04019_),
    .B1(_03878_),
    .Y(_04021_));
 sky130_fd_sc_hd__a211oi_1 _09893_ (.A1(_03920_),
    .A2(_03922_),
    .B1(_04020_),
    .C1(_04021_),
    .Y(_04022_));
 sky130_fd_sc_hd__o211a_1 _09894_ (.A1(_04020_),
    .A2(_04021_),
    .B1(_03920_),
    .C1(_03922_),
    .X(_04023_));
 sky130_fd_sc_hd__or3_2 _09895_ (.A(_03982_),
    .B(_04022_),
    .C(_04023_),
    .X(_04024_));
 sky130_fd_sc_hd__o21ai_1 _09896_ (.A1(_04022_),
    .A2(_04023_),
    .B1(_03982_),
    .Y(_04025_));
 sky130_fd_sc_hd__o211a_1 _09897_ (.A1(_03883_),
    .A2(_03928_),
    .B1(_04024_),
    .C1(_04025_),
    .X(_04026_));
 sky130_fd_sc_hd__a211oi_1 _09898_ (.A1(_04024_),
    .A2(_04025_),
    .B1(_03883_),
    .C1(_03928_),
    .Y(_04028_));
 sky130_fd_sc_hd__a211oi_2 _09899_ (.A1(_03924_),
    .A2(_03926_),
    .B1(_04026_),
    .C1(_04028_),
    .Y(_04029_));
 sky130_fd_sc_hd__o211a_1 _09900_ (.A1(_04026_),
    .A2(_04028_),
    .B1(_03924_),
    .C1(_03926_),
    .X(_04030_));
 sky130_fd_sc_hd__a211oi_2 _09901_ (.A1(_03933_),
    .A2(_03935_),
    .B1(_04029_),
    .C1(_04030_),
    .Y(_04031_));
 sky130_fd_sc_hd__o211a_1 _09902_ (.A1(_04029_),
    .A2(_04030_),
    .B1(_03933_),
    .C1(_03935_),
    .X(_04032_));
 sky130_fd_sc_hd__a211oi_2 _09903_ (.A1(_03896_),
    .A2(_03900_),
    .B1(_04031_),
    .C1(_04032_),
    .Y(_04033_));
 sky130_fd_sc_hd__o211a_1 _09904_ (.A1(_04031_),
    .A2(_04032_),
    .B1(_03896_),
    .C1(_03900_),
    .X(_04034_));
 sky130_fd_sc_hd__o211a_1 _09905_ (.A1(_04033_),
    .A2(_04034_),
    .B1(_03938_),
    .C1(_03942_),
    .X(_04035_));
 sky130_fd_sc_hd__a211oi_1 _09906_ (.A1(_03938_),
    .A2(_03942_),
    .B1(_04033_),
    .C1(_04034_),
    .Y(_04036_));
 sky130_fd_sc_hd__nor2_1 _09907_ (.A(_04035_),
    .B(_04036_),
    .Y(_04037_));
 sky130_fd_sc_hd__a21oi_1 _09908_ (.A1(_03947_),
    .A2(_03950_),
    .B1(_03946_),
    .Y(_04039_));
 sky130_fd_sc_hd__xnor2_1 _09909_ (.A(_04037_),
    .B(_04039_),
    .Y(net106));
 sky130_fd_sc_hd__nor2_1 _09910_ (.A(_03742_),
    .B(_03953_),
    .Y(_04040_));
 sky130_fd_sc_hd__xor2_1 _09911_ (.A(_03956_),
    .B(_04040_),
    .X(_04041_));
 sky130_fd_sc_hd__and4_1 _09912_ (.A(net329),
    .B(net321),
    .C(net554),
    .D(net540),
    .X(_04042_));
 sky130_fd_sc_hd__a22o_1 _09913_ (.A1(net321),
    .A2(net556),
    .B1(net540),
    .B2(net329),
    .X(_04043_));
 sky130_fd_sc_hd__and2b_1 _09914_ (.A_N(_04042_),
    .B(_04043_),
    .X(_04044_));
 sky130_fd_sc_hd__nand2_1 _09915_ (.A(net314),
    .B(net561),
    .Y(_04045_));
 sky130_fd_sc_hd__xnor2_1 _09916_ (.A(_04044_),
    .B(_04045_),
    .Y(_04046_));
 sky130_fd_sc_hd__nand2_1 _09917_ (.A(net352),
    .B(net512),
    .Y(_04047_));
 sky130_fd_sc_hd__nand4_1 _09918_ (.A(net359),
    .B(net351),
    .C(net526),
    .D(net512),
    .Y(_04049_));
 sky130_fd_sc_hd__a22o_1 _09919_ (.A1(net351),
    .A2(net526),
    .B1(net512),
    .B2(net359),
    .X(_04050_));
 sky130_fd_sc_hd__a22o_1 _09920_ (.A1(net336),
    .A2(net534),
    .B1(_04049_),
    .B2(_04050_),
    .X(_04051_));
 sky130_fd_sc_hd__nand4_1 _09921_ (.A(net336),
    .B(net534),
    .C(_04049_),
    .D(_04050_),
    .Y(_04052_));
 sky130_fd_sc_hd__nand2_1 _09922_ (.A(_03967_),
    .B(_03970_),
    .Y(_04053_));
 sky130_fd_sc_hd__and3_1 _09923_ (.A(_04051_),
    .B(_04052_),
    .C(_04053_),
    .X(_04054_));
 sky130_fd_sc_hd__a21o_1 _09924_ (.A1(_04051_),
    .A2(_04052_),
    .B1(_04053_),
    .X(_04055_));
 sky130_fd_sc_hd__and2b_1 _09925_ (.A_N(_04054_),
    .B(_04055_),
    .X(_04056_));
 sky130_fd_sc_hd__xnor2_1 _09926_ (.A(_04046_),
    .B(_04056_),
    .Y(_04057_));
 sky130_fd_sc_hd__and2_1 _09927_ (.A(_04041_),
    .B(_04057_),
    .X(_04058_));
 sky130_fd_sc_hd__nor2_1 _09928_ (.A(_04041_),
    .B(_04057_),
    .Y(_04060_));
 sky130_fd_sc_hd__a211o_1 _09929_ (.A1(_03959_),
    .A2(_03978_),
    .B1(_04058_),
    .C1(_04060_),
    .X(_04061_));
 sky130_fd_sc_hd__o211ai_1 _09930_ (.A1(_04058_),
    .A2(_04060_),
    .B1(_03959_),
    .C1(_03978_),
    .Y(_04062_));
 sky130_fd_sc_hd__nand2_1 _09931_ (.A(_04015_),
    .B(_04018_),
    .Y(_04063_));
 sky130_fd_sc_hd__and4_1 _09932_ (.A(net592),
    .B(net585),
    .C(net277),
    .D(net269),
    .X(_04064_));
 sky130_fd_sc_hd__a22oi_1 _09933_ (.A1(net585),
    .A2(net277),
    .B1(net269),
    .B2(net592),
    .Y(_04065_));
 sky130_fd_sc_hd__o2bb2a_1 _09934_ (.A1_N(net609),
    .A2_N(net261),
    .B1(_04064_),
    .B2(_04065_),
    .X(_04066_));
 sky130_fd_sc_hd__and4bb_1 _09935_ (.A_N(_04064_),
    .B_N(_04065_),
    .C(net609),
    .D(net261),
    .X(_04067_));
 sky130_fd_sc_hd__nor2_1 _09936_ (.A(_04066_),
    .B(_04067_),
    .Y(_04068_));
 sky130_fd_sc_hd__nor2_1 _09937_ (.A(_03983_),
    .B(_03986_),
    .Y(_04069_));
 sky130_fd_sc_hd__xnor2_1 _09938_ (.A(_04068_),
    .B(_04069_),
    .Y(_04071_));
 sky130_fd_sc_hd__nand2_1 _09939_ (.A(net617),
    .B(net250),
    .Y(_04072_));
 sky130_fd_sc_hd__inv_2 _09940_ (.A(_04072_),
    .Y(_04073_));
 sky130_fd_sc_hd__nand2_1 _09941_ (.A(_04071_),
    .B(_04073_),
    .Y(_04074_));
 sky130_fd_sc_hd__xnor2_1 _09942_ (.A(_04071_),
    .B(_04073_),
    .Y(_04075_));
 sky130_fd_sc_hd__a21oi_1 _09943_ (.A1(_03990_),
    .A2(_03991_),
    .B1(_03989_),
    .Y(_04076_));
 sky130_fd_sc_hd__xor2_1 _09944_ (.A(_04075_),
    .B(_04076_),
    .X(_04077_));
 sky130_fd_sc_hd__a21oi_1 _09945_ (.A1(net166),
    .A2(net244),
    .B1(_04077_),
    .Y(_04078_));
 sky130_fd_sc_hd__and3_1 _09946_ (.A(net166),
    .B(net244),
    .C(_04077_),
    .X(_04079_));
 sky130_fd_sc_hd__nor2_1 _09947_ (.A(_04078_),
    .B(_04079_),
    .Y(_04080_));
 sky130_fd_sc_hd__a21o_1 _09948_ (.A1(_03966_),
    .A2(_03974_),
    .B1(_03972_),
    .X(_04082_));
 sky130_fd_sc_hd__nand2_1 _09949_ (.A(_04002_),
    .B(_04006_),
    .Y(_04083_));
 sky130_fd_sc_hd__a31o_1 _09950_ (.A1(net314),
    .A2(net569),
    .A3(_03963_),
    .B1(_03961_),
    .X(_04084_));
 sky130_fd_sc_hd__nand4_2 _09951_ (.A(net576),
    .B(net569),
    .C(net307),
    .D(net292),
    .Y(_04085_));
 sky130_fd_sc_hd__a22o_1 _09952_ (.A1(net569),
    .A2(net307),
    .B1(net292),
    .B2(net576),
    .X(_04086_));
 sky130_fd_sc_hd__a22o_1 _09953_ (.A1(net582),
    .A2(net285),
    .B1(_04085_),
    .B2(_04086_),
    .X(_04087_));
 sky130_fd_sc_hd__nand4_2 _09954_ (.A(net582),
    .B(net285),
    .C(_04085_),
    .D(_04086_),
    .Y(_04088_));
 sky130_fd_sc_hd__nand3_2 _09955_ (.A(_04084_),
    .B(_04087_),
    .C(_04088_),
    .Y(_04089_));
 sky130_fd_sc_hd__a21o_1 _09956_ (.A1(_04087_),
    .A2(_04088_),
    .B1(_04084_),
    .X(_04090_));
 sky130_fd_sc_hd__nand3_2 _09957_ (.A(_04083_),
    .B(_04089_),
    .C(_04090_),
    .Y(_04091_));
 sky130_fd_sc_hd__a21o_1 _09958_ (.A1(_04089_),
    .A2(_04090_),
    .B1(_04083_),
    .X(_04093_));
 sky130_fd_sc_hd__and3_2 _09959_ (.A(_04082_),
    .B(_04091_),
    .C(_04093_),
    .X(_04094_));
 sky130_fd_sc_hd__a21oi_1 _09960_ (.A1(_04091_),
    .A2(_04093_),
    .B1(_04082_),
    .Y(_04095_));
 sky130_fd_sc_hd__a211oi_1 _09961_ (.A1(_04007_),
    .A2(_04009_),
    .B1(_04094_),
    .C1(_04095_),
    .Y(_04096_));
 sky130_fd_sc_hd__a211o_1 _09962_ (.A1(_04007_),
    .A2(_04009_),
    .B1(_04094_),
    .C1(_04095_),
    .X(_04097_));
 sky130_fd_sc_hd__o211ai_2 _09963_ (.A1(_04094_),
    .A2(_04095_),
    .B1(_04007_),
    .C1(_04009_),
    .Y(_04098_));
 sky130_fd_sc_hd__o211ai_2 _09964_ (.A1(_04011_),
    .A2(_04013_),
    .B1(_04097_),
    .C1(_04098_),
    .Y(_04099_));
 sky130_fd_sc_hd__a211o_1 _09965_ (.A1(_04097_),
    .A2(_04098_),
    .B1(_04011_),
    .C1(_04013_),
    .X(_04100_));
 sky130_fd_sc_hd__nand3_1 _09966_ (.A(_04080_),
    .B(_04099_),
    .C(_04100_),
    .Y(_04101_));
 sky130_fd_sc_hd__a21o_1 _09967_ (.A1(_04099_),
    .A2(_04100_),
    .B1(_04080_),
    .X(_04102_));
 sky130_fd_sc_hd__nand3_2 _09968_ (.A(_03980_),
    .B(_04101_),
    .C(_04102_),
    .Y(_04104_));
 sky130_fd_sc_hd__a21o_1 _09969_ (.A1(_04101_),
    .A2(_04102_),
    .B1(_03980_),
    .X(_04105_));
 sky130_fd_sc_hd__nand3_1 _09970_ (.A(_04063_),
    .B(_04104_),
    .C(_04105_),
    .Y(_04106_));
 sky130_fd_sc_hd__a21o_1 _09971_ (.A1(_04104_),
    .A2(_04105_),
    .B1(_04063_),
    .X(_04107_));
 sky130_fd_sc_hd__and4_1 _09972_ (.A(_04061_),
    .B(_04062_),
    .C(_04106_),
    .D(_04107_),
    .X(_04108_));
 sky130_fd_sc_hd__a22oi_1 _09973_ (.A1(_04061_),
    .A2(_04062_),
    .B1(_04106_),
    .B2(_04107_),
    .Y(_04109_));
 sky130_fd_sc_hd__or3_1 _09974_ (.A(_04024_),
    .B(_04108_),
    .C(_04109_),
    .X(_04110_));
 sky130_fd_sc_hd__o21ai_1 _09975_ (.A1(_04108_),
    .A2(_04109_),
    .B1(_04024_),
    .Y(_04111_));
 sky130_fd_sc_hd__nand2_1 _09976_ (.A(_04110_),
    .B(_04111_),
    .Y(_04112_));
 sky130_fd_sc_hd__nor2_1 _09977_ (.A(_04020_),
    .B(_04022_),
    .Y(_04113_));
 sky130_fd_sc_hd__or2_1 _09978_ (.A(_04112_),
    .B(_04113_),
    .X(_04115_));
 sky130_fd_sc_hd__xor2_1 _09979_ (.A(_04112_),
    .B(_04113_),
    .X(_04116_));
 sky130_fd_sc_hd__nor2_1 _09980_ (.A(_04026_),
    .B(_04029_),
    .Y(_04117_));
 sky130_fd_sc_hd__and2b_1 _09981_ (.A_N(_04117_),
    .B(_04116_),
    .X(_04118_));
 sky130_fd_sc_hd__xnor2_1 _09982_ (.A(_04116_),
    .B(_04117_),
    .Y(_04119_));
 sky130_fd_sc_hd__o21a_1 _09983_ (.A1(_03992_),
    .A2(_03993_),
    .B1(_03997_),
    .X(_04120_));
 sky130_fd_sc_hd__and2b_1 _09984_ (.A_N(_04120_),
    .B(_04119_),
    .X(_04121_));
 sky130_fd_sc_hd__and2b_1 _09985_ (.A_N(_04119_),
    .B(_04120_),
    .X(_04122_));
 sky130_fd_sc_hd__or2_1 _09986_ (.A(_04121_),
    .B(_04122_),
    .X(_04123_));
 sky130_fd_sc_hd__nor2_1 _09987_ (.A(_04031_),
    .B(_04033_),
    .Y(_04124_));
 sky130_fd_sc_hd__nor2_1 _09988_ (.A(_04123_),
    .B(_04124_),
    .Y(_04126_));
 sky130_fd_sc_hd__and2_1 _09989_ (.A(_04123_),
    .B(_04124_),
    .X(_04127_));
 sky130_fd_sc_hd__nor2_1 _09990_ (.A(_04126_),
    .B(_04127_),
    .Y(_04128_));
 sky130_fd_sc_hd__a31oi_1 _09991_ (.A1(_03508_),
    .A2(_03509_),
    .A3(_03621_),
    .B1(_03737_),
    .Y(_04129_));
 sky130_fd_sc_hd__nand2_1 _09992_ (.A(_03947_),
    .B(_04037_),
    .Y(_04130_));
 sky130_fd_sc_hd__or2_1 _09993_ (.A(_03949_),
    .B(_04130_),
    .X(_04131_));
 sky130_fd_sc_hd__nor2_1 _09994_ (.A(_03946_),
    .B(_04036_),
    .Y(_04132_));
 sky130_fd_sc_hd__o22a_1 _09995_ (.A1(_03948_),
    .A2(_04130_),
    .B1(_04132_),
    .B2(_04035_),
    .X(_04133_));
 sky130_fd_sc_hd__o21a_2 _09996_ (.A1(_04129_),
    .A2(_04131_),
    .B1(_04133_),
    .X(_04134_));
 sky130_fd_sc_hd__or4_4 _09997_ (.A(_03259_),
    .B(_03392_),
    .C(_03738_),
    .D(_04131_),
    .X(_04135_));
 sky130_fd_sc_hd__and2_1 _09998_ (.A(_03265_),
    .B(_04134_),
    .X(_04137_));
 sky130_fd_sc_hd__a22oi_4 _09999_ (.A1(_04134_),
    .A2(_04135_),
    .B1(_04137_),
    .B2(_03267_),
    .Y(_04138_));
 sky130_fd_sc_hd__a22o_1 _10000_ (.A1(_04134_),
    .A2(_04135_),
    .B1(_04137_),
    .B2(_03267_),
    .X(_04139_));
 sky130_fd_sc_hd__xnor2_1 _10001_ (.A(_04128_),
    .B(_04139_),
    .Y(net107));
 sky130_fd_sc_hd__and4_1 _10002_ (.A(net329),
    .B(net321),
    .C(net541),
    .D(net534),
    .X(_04140_));
 sky130_fd_sc_hd__a22o_1 _10003_ (.A1(net321),
    .A2(net541),
    .B1(net535),
    .B2(net329),
    .X(_04141_));
 sky130_fd_sc_hd__and2b_1 _10004_ (.A_N(_04140_),
    .B(_04141_),
    .X(_04142_));
 sky130_fd_sc_hd__nand2_1 _10005_ (.A(net314),
    .B(net556),
    .Y(_04143_));
 sky130_fd_sc_hd__xnor2_1 _10006_ (.A(_04142_),
    .B(_04143_),
    .Y(_04144_));
 sky130_fd_sc_hd__nand4_2 _10007_ (.A(net360),
    .B(net352),
    .C(net512),
    .D(net504),
    .Y(_04145_));
 sky130_fd_sc_hd__a22o_1 _10008_ (.A1(net352),
    .A2(net512),
    .B1(net504),
    .B2(net360),
    .X(_04147_));
 sky130_fd_sc_hd__a22o_1 _10009_ (.A1(net337),
    .A2(net526),
    .B1(_04145_),
    .B2(_04147_),
    .X(_04148_));
 sky130_fd_sc_hd__nand4_2 _10010_ (.A(net337),
    .B(net526),
    .C(_04145_),
    .D(_04147_),
    .Y(_04149_));
 sky130_fd_sc_hd__nand2_1 _10011_ (.A(_04049_),
    .B(_04052_),
    .Y(_04150_));
 sky130_fd_sc_hd__and3_1 _10012_ (.A(_04148_),
    .B(_04149_),
    .C(_04150_),
    .X(_04151_));
 sky130_fd_sc_hd__a21o_1 _10013_ (.A1(_04148_),
    .A2(_04149_),
    .B1(_04150_),
    .X(_04152_));
 sky130_fd_sc_hd__nand2b_1 _10014_ (.A_N(_04151_),
    .B(_04152_),
    .Y(_04153_));
 sky130_fd_sc_hd__xor2_1 _10015_ (.A(_04144_),
    .B(_04153_),
    .X(_04154_));
 sky130_fd_sc_hd__or3_1 _10016_ (.A(_03743_),
    .B(_03953_),
    .C(_04154_),
    .X(_04155_));
 sky130_fd_sc_hd__o21ai_1 _10017_ (.A1(_03743_),
    .A2(_03953_),
    .B1(_04154_),
    .Y(_04156_));
 sky130_fd_sc_hd__nand2_1 _10018_ (.A(_04155_),
    .B(_04156_),
    .Y(_04158_));
 sky130_fd_sc_hd__a31o_1 _10019_ (.A1(_03954_),
    .A2(_03955_),
    .A3(_04040_),
    .B1(_04060_),
    .X(_04159_));
 sky130_fd_sc_hd__and2b_1 _10020_ (.A_N(_04158_),
    .B(_04159_),
    .X(_04160_));
 sky130_fd_sc_hd__and2b_1 _10021_ (.A_N(_04159_),
    .B(_04158_),
    .X(_04161_));
 sky130_fd_sc_hd__or2_1 _10022_ (.A(_04160_),
    .B(_04161_),
    .X(_04162_));
 sky130_fd_sc_hd__nand2_1 _10023_ (.A(_04099_),
    .B(_04101_),
    .Y(_04163_));
 sky130_fd_sc_hd__and4_1 _10024_ (.A(net585),
    .B(net578),
    .C(net277),
    .D(net269),
    .X(_04164_));
 sky130_fd_sc_hd__a22oi_1 _10025_ (.A1(net578),
    .A2(net277),
    .B1(net269),
    .B2(net585),
    .Y(_04165_));
 sky130_fd_sc_hd__o2bb2a_1 _10026_ (.A1_N(net592),
    .A2_N(net261),
    .B1(_04164_),
    .B2(_04165_),
    .X(_04166_));
 sky130_fd_sc_hd__and4bb_1 _10027_ (.A_N(_04164_),
    .B_N(_04165_),
    .C(net592),
    .D(net261),
    .X(_04167_));
 sky130_fd_sc_hd__nor2_1 _10028_ (.A(_04166_),
    .B(_04167_),
    .Y(_04169_));
 sky130_fd_sc_hd__nor2_1 _10029_ (.A(_04064_),
    .B(_04067_),
    .Y(_04170_));
 sky130_fd_sc_hd__xnor2_1 _10030_ (.A(_04169_),
    .B(_04170_),
    .Y(_04171_));
 sky130_fd_sc_hd__a21o_1 _10031_ (.A1(net609),
    .A2(net250),
    .B1(_04171_),
    .X(_04172_));
 sky130_fd_sc_hd__nand3_1 _10032_ (.A(net609),
    .B(net250),
    .C(_04171_),
    .Y(_04173_));
 sky130_fd_sc_hd__nand2_1 _10033_ (.A(_04172_),
    .B(_04173_),
    .Y(_04174_));
 sky130_fd_sc_hd__o31a_1 _10034_ (.A1(_04066_),
    .A2(_04067_),
    .A3(_04069_),
    .B1(_04074_),
    .X(_04175_));
 sky130_fd_sc_hd__xnor2_1 _10035_ (.A(_04174_),
    .B(_04175_),
    .Y(_04176_));
 sky130_fd_sc_hd__nand2_1 _10036_ (.A(net617),
    .B(net244),
    .Y(_04177_));
 sky130_fd_sc_hd__or2_1 _10037_ (.A(_04176_),
    .B(_04177_),
    .X(_04178_));
 sky130_fd_sc_hd__xor2_1 _10038_ (.A(_04176_),
    .B(_04177_),
    .X(_04180_));
 sky130_fd_sc_hd__a21o_1 _10039_ (.A1(_04046_),
    .A2(_04055_),
    .B1(_04054_),
    .X(_04181_));
 sky130_fd_sc_hd__nand2_1 _10040_ (.A(_04085_),
    .B(_04088_),
    .Y(_04182_));
 sky130_fd_sc_hd__a31o_1 _10041_ (.A1(net314),
    .A2(net561),
    .A3(_04043_),
    .B1(_04042_),
    .X(_04183_));
 sky130_fd_sc_hd__nand4_2 _10042_ (.A(net569),
    .B(net307),
    .C(net561),
    .D(net292),
    .Y(_04184_));
 sky130_fd_sc_hd__a22o_1 _10043_ (.A1(net307),
    .A2(net561),
    .B1(net292),
    .B2(net569),
    .X(_04185_));
 sky130_fd_sc_hd__a22o_1 _10044_ (.A1(net576),
    .A2(net285),
    .B1(_04184_),
    .B2(_04185_),
    .X(_04186_));
 sky130_fd_sc_hd__nand4_2 _10045_ (.A(net576),
    .B(net285),
    .C(_04184_),
    .D(_04185_),
    .Y(_04187_));
 sky130_fd_sc_hd__nand3_2 _10046_ (.A(_04183_),
    .B(_04186_),
    .C(_04187_),
    .Y(_04188_));
 sky130_fd_sc_hd__a21o_1 _10047_ (.A1(_04186_),
    .A2(_04187_),
    .B1(_04183_),
    .X(_04189_));
 sky130_fd_sc_hd__nand3_2 _10048_ (.A(_04182_),
    .B(_04188_),
    .C(_04189_),
    .Y(_04191_));
 sky130_fd_sc_hd__a21o_1 _10049_ (.A1(_04188_),
    .A2(_04189_),
    .B1(_04182_),
    .X(_04192_));
 sky130_fd_sc_hd__and3_2 _10050_ (.A(_04181_),
    .B(_04191_),
    .C(_04192_),
    .X(_04193_));
 sky130_fd_sc_hd__a21oi_2 _10051_ (.A1(_04191_),
    .A2(_04192_),
    .B1(_04181_),
    .Y(_04194_));
 sky130_fd_sc_hd__a211oi_2 _10052_ (.A1(_04089_),
    .A2(_04091_),
    .B1(_04193_),
    .C1(_04194_),
    .Y(_04195_));
 sky130_fd_sc_hd__a211o_1 _10053_ (.A1(_04089_),
    .A2(_04091_),
    .B1(_04193_),
    .C1(_04194_),
    .X(_04196_));
 sky130_fd_sc_hd__o211ai_2 _10054_ (.A1(_04193_),
    .A2(_04194_),
    .B1(_04089_),
    .C1(_04091_),
    .Y(_04197_));
 sky130_fd_sc_hd__o211a_1 _10055_ (.A1(_04094_),
    .A2(_04096_),
    .B1(_04196_),
    .C1(_04197_),
    .X(_04198_));
 sky130_fd_sc_hd__o211ai_1 _10056_ (.A1(_04094_),
    .A2(_04096_),
    .B1(_04196_),
    .C1(_04197_),
    .Y(_04199_));
 sky130_fd_sc_hd__a211o_1 _10057_ (.A1(_04196_),
    .A2(_04197_),
    .B1(_04094_),
    .C1(_04096_),
    .X(_04200_));
 sky130_fd_sc_hd__and3_1 _10058_ (.A(_04180_),
    .B(_04199_),
    .C(_04200_),
    .X(_04202_));
 sky130_fd_sc_hd__a21oi_1 _10059_ (.A1(_04199_),
    .A2(_04200_),
    .B1(_04180_),
    .Y(_04203_));
 sky130_fd_sc_hd__nor3_1 _10060_ (.A(_04061_),
    .B(_04202_),
    .C(_04203_),
    .Y(_04204_));
 sky130_fd_sc_hd__or3_1 _10061_ (.A(_04061_),
    .B(_04202_),
    .C(_04203_),
    .X(_04205_));
 sky130_fd_sc_hd__o21ai_1 _10062_ (.A1(_04202_),
    .A2(_04203_),
    .B1(_04061_),
    .Y(_04206_));
 sky130_fd_sc_hd__and3_1 _10063_ (.A(_04163_),
    .B(_04205_),
    .C(_04206_),
    .X(_04207_));
 sky130_fd_sc_hd__a21oi_1 _10064_ (.A1(_04205_),
    .A2(_04206_),
    .B1(_04163_),
    .Y(_04208_));
 sky130_fd_sc_hd__or3_1 _10065_ (.A(_04162_),
    .B(_04207_),
    .C(_04208_),
    .X(_04209_));
 sky130_fd_sc_hd__o21ai_1 _10066_ (.A1(_04207_),
    .A2(_04208_),
    .B1(_04162_),
    .Y(_04210_));
 sky130_fd_sc_hd__and3_1 _10067_ (.A(_04108_),
    .B(_04209_),
    .C(_04210_),
    .X(_04211_));
 sky130_fd_sc_hd__a21oi_1 _10068_ (.A1(_04209_),
    .A2(_04210_),
    .B1(_04108_),
    .Y(_04213_));
 sky130_fd_sc_hd__a211oi_2 _10069_ (.A1(_04104_),
    .A2(_04106_),
    .B1(_04211_),
    .C1(_04213_),
    .Y(_04214_));
 sky130_fd_sc_hd__o211a_1 _10070_ (.A1(_04211_),
    .A2(_04213_),
    .B1(_04104_),
    .C1(_04106_),
    .X(_04215_));
 sky130_fd_sc_hd__a211oi_1 _10071_ (.A1(_04110_),
    .A2(_04115_),
    .B1(_04214_),
    .C1(_04215_),
    .Y(_04216_));
 sky130_fd_sc_hd__o211a_1 _10072_ (.A1(_04214_),
    .A2(_04215_),
    .B1(_04110_),
    .C1(_04115_),
    .X(_04217_));
 sky130_fd_sc_hd__nor2_1 _10073_ (.A(_04216_),
    .B(_04217_),
    .Y(_04218_));
 sky130_fd_sc_hd__o21ba_1 _10074_ (.A1(_04075_),
    .A2(_04076_),
    .B1_N(_04079_),
    .X(_04219_));
 sky130_fd_sc_hd__xnor2_1 _10075_ (.A(_04218_),
    .B(_04219_),
    .Y(_04220_));
 sky130_fd_sc_hd__nor3_1 _10076_ (.A(_04118_),
    .B(_04121_),
    .C(_04220_),
    .Y(_04221_));
 sky130_fd_sc_hd__or3_1 _10077_ (.A(_04118_),
    .B(_04121_),
    .C(_04220_),
    .X(_04222_));
 sky130_fd_sc_hd__o21a_1 _10078_ (.A1(_04118_),
    .A2(_04121_),
    .B1(_04220_),
    .X(_04224_));
 sky130_fd_sc_hd__nor2_1 _10079_ (.A(_04221_),
    .B(_04224_),
    .Y(_04225_));
 sky130_fd_sc_hd__a21oi_1 _10080_ (.A1(_04128_),
    .A2(_04138_),
    .B1(_04126_),
    .Y(_04226_));
 sky130_fd_sc_hd__xnor2_1 _10081_ (.A(_04225_),
    .B(_04226_),
    .Y(net108));
 sky130_fd_sc_hd__nand2_1 _10082_ (.A(net337),
    .B(net505),
    .Y(_04227_));
 sky130_fd_sc_hd__a22o_1 _10083_ (.A1(net337),
    .A2(net512),
    .B1(net505),
    .B2(net352),
    .X(_04228_));
 sky130_fd_sc_hd__o21a_1 _10084_ (.A1(_04047_),
    .A2(_04227_),
    .B1(_04228_),
    .X(_04229_));
 sky130_fd_sc_hd__o21ai_1 _10085_ (.A1(_04047_),
    .A2(_04227_),
    .B1(_04228_),
    .Y(_04230_));
 sky130_fd_sc_hd__nand3_1 _10086_ (.A(_04145_),
    .B(_04149_),
    .C(_04230_),
    .Y(_04231_));
 sky130_fd_sc_hd__inv_2 _10087_ (.A(_04231_),
    .Y(_04232_));
 sky130_fd_sc_hd__a21boi_1 _10088_ (.A1(_04145_),
    .A2(_04149_),
    .B1_N(_04229_),
    .Y(_04234_));
 sky130_fd_sc_hd__nor2_1 _10089_ (.A(_04232_),
    .B(_04234_),
    .Y(_04235_));
 sky130_fd_sc_hd__and4_1 _10090_ (.A(net329),
    .B(net321),
    .C(net535),
    .D(net526),
    .X(_04236_));
 sky130_fd_sc_hd__a22o_1 _10091_ (.A1(net321),
    .A2(net535),
    .B1(net527),
    .B2(net329),
    .X(_04237_));
 sky130_fd_sc_hd__and2b_1 _10092_ (.A_N(_04236_),
    .B(_04237_),
    .X(_04238_));
 sky130_fd_sc_hd__nand2_1 _10093_ (.A(net315),
    .B(net541),
    .Y(_04239_));
 sky130_fd_sc_hd__xnor2_1 _10094_ (.A(_04238_),
    .B(_04239_),
    .Y(_04240_));
 sky130_fd_sc_hd__xnor2_1 _10095_ (.A(_04235_),
    .B(_04240_),
    .Y(_04241_));
 sky130_fd_sc_hd__or2_1 _10096_ (.A(_04155_),
    .B(_04241_),
    .X(_04242_));
 sky130_fd_sc_hd__nand2_1 _10097_ (.A(_04155_),
    .B(_04241_),
    .Y(_04243_));
 sky130_fd_sc_hd__nand2_1 _10098_ (.A(_04242_),
    .B(_04243_),
    .Y(_04245_));
 sky130_fd_sc_hd__and4_1 _10099_ (.A(net578),
    .B(net572),
    .C(net278),
    .D(net270),
    .X(_04246_));
 sky130_fd_sc_hd__a22oi_1 _10100_ (.A1(net572),
    .A2(net278),
    .B1(net270),
    .B2(net578),
    .Y(_04247_));
 sky130_fd_sc_hd__nor2_1 _10101_ (.A(_04246_),
    .B(_04247_),
    .Y(_04248_));
 sky130_fd_sc_hd__nand2_1 _10102_ (.A(net585),
    .B(net262),
    .Y(_04249_));
 sky130_fd_sc_hd__xnor2_1 _10103_ (.A(_04248_),
    .B(_04249_),
    .Y(_04250_));
 sky130_fd_sc_hd__nor3_1 _10104_ (.A(_04164_),
    .B(_04167_),
    .C(_04250_),
    .Y(_04251_));
 sky130_fd_sc_hd__o21a_1 _10105_ (.A1(_04164_),
    .A2(_04167_),
    .B1(_04250_),
    .X(_04252_));
 sky130_fd_sc_hd__nor2_1 _10106_ (.A(_04251_),
    .B(_04252_),
    .Y(_04253_));
 sky130_fd_sc_hd__nand2_1 _10107_ (.A(net592),
    .B(net250),
    .Y(_04254_));
 sky130_fd_sc_hd__xor2_1 _10108_ (.A(_04253_),
    .B(_04254_),
    .X(_04256_));
 sky130_fd_sc_hd__o31a_1 _10109_ (.A1(_04166_),
    .A2(_04167_),
    .A3(_04170_),
    .B1(_04173_),
    .X(_04257_));
 sky130_fd_sc_hd__or2_1 _10110_ (.A(_04256_),
    .B(_04257_),
    .X(_04258_));
 sky130_fd_sc_hd__xnor2_1 _10111_ (.A(_04256_),
    .B(_04257_),
    .Y(_04259_));
 sky130_fd_sc_hd__nand2_1 _10112_ (.A(net609),
    .B(net244),
    .Y(_04260_));
 sky130_fd_sc_hd__or2_1 _10113_ (.A(_04259_),
    .B(_04260_),
    .X(_04261_));
 sky130_fd_sc_hd__xor2_1 _10114_ (.A(_04259_),
    .B(_04260_),
    .X(_04262_));
 sky130_fd_sc_hd__a21o_1 _10115_ (.A1(_04144_),
    .A2(_04152_),
    .B1(_04151_),
    .X(_04263_));
 sky130_fd_sc_hd__nand2_1 _10116_ (.A(_04184_),
    .B(_04187_),
    .Y(_04264_));
 sky130_fd_sc_hd__a31o_1 _10117_ (.A1(net315),
    .A2(net556),
    .A3(_04141_),
    .B1(_04140_),
    .X(_04265_));
 sky130_fd_sc_hd__nand4_2 _10118_ (.A(net307),
    .B(net561),
    .C(net293),
    .D(net555),
    .Y(_04267_));
 sky130_fd_sc_hd__a22o_1 _10119_ (.A1(net561),
    .A2(net293),
    .B1(net555),
    .B2(net307),
    .X(_04268_));
 sky130_fd_sc_hd__a22o_1 _10120_ (.A1(net569),
    .A2(net286),
    .B1(_04267_),
    .B2(_04268_),
    .X(_04269_));
 sky130_fd_sc_hd__nand4_2 _10121_ (.A(net569),
    .B(net286),
    .C(_04267_),
    .D(_04268_),
    .Y(_04270_));
 sky130_fd_sc_hd__nand3_2 _10122_ (.A(_04265_),
    .B(_04269_),
    .C(_04270_),
    .Y(_04271_));
 sky130_fd_sc_hd__a21o_1 _10123_ (.A1(_04269_),
    .A2(_04270_),
    .B1(_04265_),
    .X(_04272_));
 sky130_fd_sc_hd__nand3_1 _10124_ (.A(_04264_),
    .B(_04271_),
    .C(_04272_),
    .Y(_04273_));
 sky130_fd_sc_hd__a21o_1 _10125_ (.A1(_04271_),
    .A2(_04272_),
    .B1(_04264_),
    .X(_04274_));
 sky130_fd_sc_hd__and3_2 _10126_ (.A(_04263_),
    .B(_04273_),
    .C(_04274_),
    .X(_04275_));
 sky130_fd_sc_hd__a21oi_1 _10127_ (.A1(_04273_),
    .A2(_04274_),
    .B1(_04263_),
    .Y(_04276_));
 sky130_fd_sc_hd__a211oi_1 _10128_ (.A1(_04188_),
    .A2(_04191_),
    .B1(_04275_),
    .C1(_04276_),
    .Y(_04278_));
 sky130_fd_sc_hd__a211o_1 _10129_ (.A1(_04188_),
    .A2(_04191_),
    .B1(_04275_),
    .C1(_04276_),
    .X(_04279_));
 sky130_fd_sc_hd__o211ai_2 _10130_ (.A1(_04275_),
    .A2(_04276_),
    .B1(_04188_),
    .C1(_04191_),
    .Y(_04280_));
 sky130_fd_sc_hd__o211ai_4 _10131_ (.A1(_04193_),
    .A2(_04195_),
    .B1(_04279_),
    .C1(_04280_),
    .Y(_04281_));
 sky130_fd_sc_hd__a211o_1 _10132_ (.A1(_04279_),
    .A2(_04280_),
    .B1(_04193_),
    .C1(_04195_),
    .X(_04282_));
 sky130_fd_sc_hd__nand3_2 _10133_ (.A(_04262_),
    .B(_04281_),
    .C(_04282_),
    .Y(_04283_));
 sky130_fd_sc_hd__a21o_1 _10134_ (.A1(_04281_),
    .A2(_04282_),
    .B1(_04262_),
    .X(_04284_));
 sky130_fd_sc_hd__nand3_2 _10135_ (.A(_04160_),
    .B(_04283_),
    .C(_04284_),
    .Y(_04285_));
 sky130_fd_sc_hd__a21o_1 _10136_ (.A1(_04283_),
    .A2(_04284_),
    .B1(_04160_),
    .X(_04286_));
 sky130_fd_sc_hd__o211a_1 _10137_ (.A1(_04198_),
    .A2(_04202_),
    .B1(_04285_),
    .C1(_04286_),
    .X(_04287_));
 sky130_fd_sc_hd__inv_2 _10138_ (.A(_04287_),
    .Y(_04289_));
 sky130_fd_sc_hd__a211oi_1 _10139_ (.A1(_04285_),
    .A2(_04286_),
    .B1(_04198_),
    .C1(_04202_),
    .Y(_04290_));
 sky130_fd_sc_hd__nor3_1 _10140_ (.A(_04245_),
    .B(_04287_),
    .C(_04290_),
    .Y(_04291_));
 sky130_fd_sc_hd__o21a_1 _10141_ (.A1(_04287_),
    .A2(_04290_),
    .B1(_04245_),
    .X(_04292_));
 sky130_fd_sc_hd__or3_2 _10142_ (.A(_04209_),
    .B(net131),
    .C(_04292_),
    .X(_04293_));
 sky130_fd_sc_hd__o21ai_2 _10143_ (.A1(net131),
    .A2(_04292_),
    .B1(_04209_),
    .Y(_04294_));
 sky130_fd_sc_hd__o211ai_4 _10144_ (.A1(net137),
    .A2(_04207_),
    .B1(_04293_),
    .C1(_04294_),
    .Y(_04295_));
 sky130_fd_sc_hd__a211o_1 _10145_ (.A1(_04293_),
    .A2(_04294_),
    .B1(_04204_),
    .C1(_04207_),
    .X(_04296_));
 sky130_fd_sc_hd__o211ai_2 _10146_ (.A1(_04211_),
    .A2(_04214_),
    .B1(_04295_),
    .C1(_04296_),
    .Y(_04297_));
 sky130_fd_sc_hd__a211o_1 _10147_ (.A1(_04295_),
    .A2(_04296_),
    .B1(_04211_),
    .C1(_04214_),
    .X(_04298_));
 sky130_fd_sc_hd__o21a_1 _10148_ (.A1(_04174_),
    .A2(_04175_),
    .B1(_04178_),
    .X(_04300_));
 sky130_fd_sc_hd__inv_2 _10149_ (.A(_04300_),
    .Y(_04301_));
 sky130_fd_sc_hd__nand3_1 _10150_ (.A(_04297_),
    .B(_04298_),
    .C(_04301_),
    .Y(_04302_));
 sky130_fd_sc_hd__a21o_1 _10151_ (.A1(_04297_),
    .A2(_04298_),
    .B1(_04301_),
    .X(_04303_));
 sky130_fd_sc_hd__nand2_1 _10152_ (.A(_04302_),
    .B(_04303_),
    .Y(_04304_));
 sky130_fd_sc_hd__o21ba_1 _10153_ (.A1(_04217_),
    .A2(_04219_),
    .B1_N(_04216_),
    .X(_04305_));
 sky130_fd_sc_hd__nor2_1 _10154_ (.A(_04304_),
    .B(_04305_),
    .Y(_04306_));
 sky130_fd_sc_hd__nand2_1 _10155_ (.A(_04304_),
    .B(_04305_),
    .Y(_04307_));
 sky130_fd_sc_hd__nand2b_1 _10156_ (.A_N(_04306_),
    .B(_04307_),
    .Y(_04308_));
 sky130_fd_sc_hd__a21oi_1 _10157_ (.A1(_04126_),
    .A2(_04222_),
    .B1(_04224_),
    .Y(_04309_));
 sky130_fd_sc_hd__nand2_1 _10158_ (.A(_04128_),
    .B(_04225_),
    .Y(_04311_));
 sky130_fd_sc_hd__o21ai_1 _10159_ (.A1(_04139_),
    .A2(_04311_),
    .B1(_04309_),
    .Y(_04312_));
 sky130_fd_sc_hd__xnor2_1 _10160_ (.A(_04308_),
    .B(_04312_),
    .Y(net110));
 sky130_fd_sc_hd__and3_1 _10161_ (.A(net337),
    .B(net505),
    .C(_04047_),
    .X(_04313_));
 sky130_fd_sc_hd__and4_1 _10162_ (.A(net334),
    .B(net322),
    .C(net527),
    .D(net511),
    .X(_04314_));
 sky130_fd_sc_hd__a22oi_1 _10163_ (.A1(net322),
    .A2(net527),
    .B1(net511),
    .B2(net334),
    .Y(_04315_));
 sky130_fd_sc_hd__nor2_1 _10164_ (.A(_04314_),
    .B(_04315_),
    .Y(_04316_));
 sky130_fd_sc_hd__nand2_1 _10165_ (.A(net315),
    .B(net535),
    .Y(_04317_));
 sky130_fd_sc_hd__xnor2_1 _10166_ (.A(_04316_),
    .B(_04317_),
    .Y(_04318_));
 sky130_fd_sc_hd__inv_2 _10167_ (.A(_04318_),
    .Y(_04319_));
 sky130_fd_sc_hd__xnor2_1 _10168_ (.A(_04313_),
    .B(_04318_),
    .Y(_04321_));
 sky130_fd_sc_hd__and4_1 _10169_ (.A(net572),
    .B(net564),
    .C(net277),
    .D(net269),
    .X(_04322_));
 sky130_fd_sc_hd__a22oi_1 _10170_ (.A1(net565),
    .A2(net277),
    .B1(net269),
    .B2(net572),
    .Y(_04323_));
 sky130_fd_sc_hd__nor2_1 _10171_ (.A(_04322_),
    .B(_04323_),
    .Y(_04324_));
 sky130_fd_sc_hd__nand2_1 _10172_ (.A(net578),
    .B(net262),
    .Y(_04325_));
 sky130_fd_sc_hd__xnor2_1 _10173_ (.A(_04324_),
    .B(_04325_),
    .Y(_04326_));
 sky130_fd_sc_hd__o21ba_1 _10174_ (.A1(_04247_),
    .A2(_04249_),
    .B1_N(_04246_),
    .X(_04327_));
 sky130_fd_sc_hd__nand2b_1 _10175_ (.A_N(_04327_),
    .B(_04326_),
    .Y(_04328_));
 sky130_fd_sc_hd__xnor2_1 _10176_ (.A(_04326_),
    .B(_04327_),
    .Y(_04329_));
 sky130_fd_sc_hd__a21o_1 _10177_ (.A1(net585),
    .A2(net250),
    .B1(_04329_),
    .X(_04330_));
 sky130_fd_sc_hd__nand3_1 _10178_ (.A(net585),
    .B(net250),
    .C(_04329_),
    .Y(_04332_));
 sky130_fd_sc_hd__nand2_1 _10179_ (.A(_04330_),
    .B(_04332_),
    .Y(_04333_));
 sky130_fd_sc_hd__a31oi_2 _10180_ (.A1(net592),
    .A2(net250),
    .A3(_04253_),
    .B1(_04252_),
    .Y(_04334_));
 sky130_fd_sc_hd__or2_1 _10181_ (.A(_04333_),
    .B(_04334_),
    .X(_04335_));
 sky130_fd_sc_hd__xnor2_1 _10182_ (.A(_04333_),
    .B(_04334_),
    .Y(_04336_));
 sky130_fd_sc_hd__nand2_1 _10183_ (.A(net593),
    .B(net246),
    .Y(_04337_));
 sky130_fd_sc_hd__xor2_1 _10184_ (.A(_04336_),
    .B(_04337_),
    .X(_04338_));
 sky130_fd_sc_hd__a21o_1 _10185_ (.A1(_04231_),
    .A2(_04240_),
    .B1(_04234_),
    .X(_04339_));
 sky130_fd_sc_hd__nand2_1 _10186_ (.A(_04267_),
    .B(_04270_),
    .Y(_04340_));
 sky130_fd_sc_hd__a31o_1 _10187_ (.A1(net315),
    .A2(net541),
    .A3(_04237_),
    .B1(_04236_),
    .X(_04341_));
 sky130_fd_sc_hd__nand4_2 _10188_ (.A(net307),
    .B(net293),
    .C(net555),
    .D(net541),
    .Y(_04343_));
 sky130_fd_sc_hd__a22o_1 _10189_ (.A1(net293),
    .A2(net555),
    .B1(net541),
    .B2(net307),
    .X(_04344_));
 sky130_fd_sc_hd__a22o_1 _10190_ (.A1(net561),
    .A2(net286),
    .B1(_04343_),
    .B2(_04344_),
    .X(_04345_));
 sky130_fd_sc_hd__nand4_2 _10191_ (.A(net561),
    .B(net286),
    .C(_04343_),
    .D(_04344_),
    .Y(_04346_));
 sky130_fd_sc_hd__and3_1 _10192_ (.A(_04341_),
    .B(_04345_),
    .C(_04346_),
    .X(_04347_));
 sky130_fd_sc_hd__nand3_1 _10193_ (.A(_04341_),
    .B(_04345_),
    .C(_04346_),
    .Y(_04348_));
 sky130_fd_sc_hd__a21o_1 _10194_ (.A1(_04345_),
    .A2(_04346_),
    .B1(_04341_),
    .X(_04349_));
 sky130_fd_sc_hd__and3_1 _10195_ (.A(_04340_),
    .B(_04348_),
    .C(_04349_),
    .X(_04350_));
 sky130_fd_sc_hd__nand3_1 _10196_ (.A(_04340_),
    .B(_04348_),
    .C(_04349_),
    .Y(_04351_));
 sky130_fd_sc_hd__a21o_1 _10197_ (.A1(_04348_),
    .A2(_04349_),
    .B1(_04340_),
    .X(_04352_));
 sky130_fd_sc_hd__and3_1 _10198_ (.A(_04339_),
    .B(_04351_),
    .C(_04352_),
    .X(_04354_));
 sky130_fd_sc_hd__a21oi_1 _10199_ (.A1(_04351_),
    .A2(_04352_),
    .B1(_04339_),
    .Y(_04355_));
 sky130_fd_sc_hd__a211o_1 _10200_ (.A1(_04271_),
    .A2(_04273_),
    .B1(_04354_),
    .C1(_04355_),
    .X(_04356_));
 sky130_fd_sc_hd__o211ai_2 _10201_ (.A1(_04354_),
    .A2(_04355_),
    .B1(_04271_),
    .C1(_04273_),
    .Y(_04357_));
 sky130_fd_sc_hd__o211ai_2 _10202_ (.A1(_04275_),
    .A2(_04278_),
    .B1(_04356_),
    .C1(_04357_),
    .Y(_04358_));
 sky130_fd_sc_hd__inv_2 _10203_ (.A(_04358_),
    .Y(_04359_));
 sky130_fd_sc_hd__a211o_1 _10204_ (.A1(_04356_),
    .A2(_04357_),
    .B1(_04275_),
    .C1(_04278_),
    .X(_04360_));
 sky130_fd_sc_hd__and3_1 _10205_ (.A(_04338_),
    .B(_04358_),
    .C(_04360_),
    .X(_04361_));
 sky130_fd_sc_hd__a21oi_1 _10206_ (.A1(_04358_),
    .A2(_04360_),
    .B1(_04338_),
    .Y(_04362_));
 sky130_fd_sc_hd__nor3_1 _10207_ (.A(_04242_),
    .B(_04361_),
    .C(_04362_),
    .Y(_04363_));
 sky130_fd_sc_hd__o21a_1 _10208_ (.A1(_04361_),
    .A2(_04362_),
    .B1(_04242_),
    .X(_04365_));
 sky130_fd_sc_hd__a211oi_2 _10209_ (.A1(_04281_),
    .A2(_04283_),
    .B1(net136),
    .C1(_04365_),
    .Y(_04366_));
 sky130_fd_sc_hd__o211a_1 _10210_ (.A1(net136),
    .A2(_04365_),
    .B1(_04281_),
    .C1(_04283_),
    .X(_04367_));
 sky130_fd_sc_hd__or3_2 _10211_ (.A(_04321_),
    .B(_04366_),
    .C(_04367_),
    .X(_04368_));
 sky130_fd_sc_hd__o21ai_1 _10212_ (.A1(_04366_),
    .A2(_04367_),
    .B1(_04321_),
    .Y(_04369_));
 sky130_fd_sc_hd__and3_1 _10213_ (.A(_04291_),
    .B(_04368_),
    .C(_04369_),
    .X(_04370_));
 sky130_fd_sc_hd__a21oi_1 _10214_ (.A1(_04368_),
    .A2(_04369_),
    .B1(_04291_),
    .Y(_04371_));
 sky130_fd_sc_hd__a211oi_2 _10215_ (.A1(_04285_),
    .A2(_04289_),
    .B1(_04370_),
    .C1(_04371_),
    .Y(_04372_));
 sky130_fd_sc_hd__o211a_1 _10216_ (.A1(_04370_),
    .A2(_04371_),
    .B1(_04285_),
    .C1(_04289_),
    .X(_04373_));
 sky130_fd_sc_hd__a211oi_2 _10217_ (.A1(_04293_),
    .A2(_04295_),
    .B1(_04372_),
    .C1(_04373_),
    .Y(_04374_));
 sky130_fd_sc_hd__o211a_1 _10218_ (.A1(_04372_),
    .A2(_04373_),
    .B1(_04293_),
    .C1(_04295_),
    .X(_04376_));
 sky130_fd_sc_hd__a211oi_2 _10219_ (.A1(_04258_),
    .A2(_04261_),
    .B1(_04374_),
    .C1(_04376_),
    .Y(_04377_));
 sky130_fd_sc_hd__o211a_1 _10220_ (.A1(_04374_),
    .A2(_04376_),
    .B1(_04258_),
    .C1(_04261_),
    .X(_04378_));
 sky130_fd_sc_hd__o211a_1 _10221_ (.A1(_04377_),
    .A2(_04378_),
    .B1(_04297_),
    .C1(_04302_),
    .X(_04379_));
 sky130_fd_sc_hd__a211oi_1 _10222_ (.A1(_04297_),
    .A2(_04302_),
    .B1(_04377_),
    .C1(_04378_),
    .Y(_04380_));
 sky130_fd_sc_hd__nor2_1 _10223_ (.A(_04379_),
    .B(_04380_),
    .Y(_04381_));
 sky130_fd_sc_hd__a21oi_1 _10224_ (.A1(_04307_),
    .A2(_04312_),
    .B1(_04306_),
    .Y(_04382_));
 sky130_fd_sc_hd__xnor2_1 _10225_ (.A(_04381_),
    .B(_04382_),
    .Y(net111));
 sky130_fd_sc_hd__and4_1 _10226_ (.A(net334),
    .B(net321),
    .C(net511),
    .D(net504),
    .X(_04383_));
 sky130_fd_sc_hd__a22o_1 _10227_ (.A1(net321),
    .A2(net511),
    .B1(net504),
    .B2(net334),
    .X(_04384_));
 sky130_fd_sc_hd__and2b_1 _10228_ (.A_N(_04383_),
    .B(_04384_),
    .X(_04386_));
 sky130_fd_sc_hd__nand2_1 _10229_ (.A(net314),
    .B(net527),
    .Y(_04387_));
 sky130_fd_sc_hd__xnor2_1 _10230_ (.A(_04386_),
    .B(_04387_),
    .Y(_04388_));
 sky130_fd_sc_hd__inv_2 _10231_ (.A(_04388_),
    .Y(_04389_));
 sky130_fd_sc_hd__a21o_1 _10232_ (.A1(_04047_),
    .A2(_04319_),
    .B1(_04227_),
    .X(_04390_));
 sky130_fd_sc_hd__nand2_1 _10233_ (.A(_04343_),
    .B(_04346_),
    .Y(_04391_));
 sky130_fd_sc_hd__o21ba_1 _10234_ (.A1(_04315_),
    .A2(_04317_),
    .B1_N(_04314_),
    .X(_04392_));
 sky130_fd_sc_hd__and4_1 _10235_ (.A(net306),
    .B(net291),
    .C(net541),
    .D(net535),
    .X(_04393_));
 sky130_fd_sc_hd__a22oi_1 _10236_ (.A1(net291),
    .A2(net541),
    .B1(net535),
    .B2(net306),
    .Y(_04394_));
 sky130_fd_sc_hd__nor2_1 _10237_ (.A(_04393_),
    .B(_04394_),
    .Y(_04395_));
 sky130_fd_sc_hd__nand2_1 _10238_ (.A(net555),
    .B(net284),
    .Y(_04397_));
 sky130_fd_sc_hd__xnor2_1 _10239_ (.A(_04395_),
    .B(_04397_),
    .Y(_04398_));
 sky130_fd_sc_hd__and2b_1 _10240_ (.A_N(_04392_),
    .B(_04398_),
    .X(_04399_));
 sky130_fd_sc_hd__xnor2_1 _10241_ (.A(_04392_),
    .B(_04398_),
    .Y(_04400_));
 sky130_fd_sc_hd__xor2_1 _10242_ (.A(_04391_),
    .B(_04400_),
    .X(_04401_));
 sky130_fd_sc_hd__nand2b_1 _10243_ (.A_N(_04390_),
    .B(_04401_),
    .Y(_04402_));
 sky130_fd_sc_hd__xnor2_1 _10244_ (.A(_04390_),
    .B(_04401_),
    .Y(_04403_));
 sky130_fd_sc_hd__or3_1 _10245_ (.A(_04347_),
    .B(_04350_),
    .C(_04403_),
    .X(_04404_));
 sky130_fd_sc_hd__o21ai_1 _10246_ (.A1(_04347_),
    .A2(_04350_),
    .B1(_04403_),
    .Y(_04405_));
 sky130_fd_sc_hd__nand2b_1 _10247_ (.A_N(_04354_),
    .B(_04356_),
    .Y(_04406_));
 sky130_fd_sc_hd__a21o_1 _10248_ (.A1(_04404_),
    .A2(_04405_),
    .B1(_04406_),
    .X(_04408_));
 sky130_fd_sc_hd__nand3_1 _10249_ (.A(_04404_),
    .B(_04405_),
    .C(_04406_),
    .Y(_04409_));
 sky130_fd_sc_hd__and4_1 _10250_ (.A(net565),
    .B(net557),
    .C(net277),
    .D(net270),
    .X(_04410_));
 sky130_fd_sc_hd__a22oi_1 _10251_ (.A1(net558),
    .A2(net277),
    .B1(net270),
    .B2(net565),
    .Y(_04411_));
 sky130_fd_sc_hd__nor2_1 _10252_ (.A(_04410_),
    .B(_04411_),
    .Y(_04412_));
 sky130_fd_sc_hd__nand2_1 _10253_ (.A(net572),
    .B(net262),
    .Y(_04413_));
 sky130_fd_sc_hd__xnor2_1 _10254_ (.A(_04412_),
    .B(_04413_),
    .Y(_04414_));
 sky130_fd_sc_hd__o21ba_1 _10255_ (.A1(_04323_),
    .A2(_04325_),
    .B1_N(_04322_),
    .X(_04415_));
 sky130_fd_sc_hd__nand2b_1 _10256_ (.A_N(_04415_),
    .B(_04414_),
    .Y(_04416_));
 sky130_fd_sc_hd__xnor2_1 _10257_ (.A(_04414_),
    .B(_04415_),
    .Y(_04417_));
 sky130_fd_sc_hd__and2_1 _10258_ (.A(net583),
    .B(net251),
    .X(_04419_));
 sky130_fd_sc_hd__or2_1 _10259_ (.A(_04417_),
    .B(_04419_),
    .X(_04420_));
 sky130_fd_sc_hd__nand2_1 _10260_ (.A(_04417_),
    .B(_04419_),
    .Y(_04421_));
 sky130_fd_sc_hd__nand2_1 _10261_ (.A(_04420_),
    .B(_04421_),
    .Y(_04422_));
 sky130_fd_sc_hd__nand2_1 _10262_ (.A(_04328_),
    .B(_04332_),
    .Y(_04423_));
 sky130_fd_sc_hd__xnor2_1 _10263_ (.A(_04422_),
    .B(_04423_),
    .Y(_04424_));
 sky130_fd_sc_hd__nand2_1 _10264_ (.A(net586),
    .B(net244),
    .Y(_04425_));
 sky130_fd_sc_hd__and2_1 _10265_ (.A(net245),
    .B(_04424_),
    .X(_04426_));
 sky130_fd_sc_hd__xnor2_1 _10266_ (.A(_04424_),
    .B(_04425_),
    .Y(_04427_));
 sky130_fd_sc_hd__a21oi_1 _10267_ (.A1(_04408_),
    .A2(_04409_),
    .B1(_04427_),
    .Y(_04428_));
 sky130_fd_sc_hd__and3_1 _10268_ (.A(_04408_),
    .B(_04409_),
    .C(_04427_),
    .X(_04430_));
 sky130_fd_sc_hd__or2_1 _10269_ (.A(_04428_),
    .B(_04430_),
    .X(_04431_));
 sky130_fd_sc_hd__nor2_1 _10270_ (.A(_04359_),
    .B(_04361_),
    .Y(_04432_));
 sky130_fd_sc_hd__or2_1 _10271_ (.A(_04431_),
    .B(_04432_),
    .X(_04433_));
 sky130_fd_sc_hd__inv_2 _10272_ (.A(_04433_),
    .Y(_04434_));
 sky130_fd_sc_hd__xnor2_1 _10273_ (.A(_04431_),
    .B(_04432_),
    .Y(_04435_));
 sky130_fd_sc_hd__nor2_1 _10274_ (.A(_04389_),
    .B(_04435_),
    .Y(_04436_));
 sky130_fd_sc_hd__xnor2_1 _10275_ (.A(_04389_),
    .B(_04435_),
    .Y(_04437_));
 sky130_fd_sc_hd__xor2_1 _10276_ (.A(_04368_),
    .B(_04437_),
    .X(_04438_));
 sky130_fd_sc_hd__o21ai_1 _10277_ (.A1(_04363_),
    .A2(_04366_),
    .B1(_04438_),
    .Y(_04439_));
 sky130_fd_sc_hd__or3_1 _10278_ (.A(_04363_),
    .B(_04366_),
    .C(_04438_),
    .X(_04441_));
 sky130_fd_sc_hd__and2_1 _10279_ (.A(_04439_),
    .B(_04441_),
    .X(_04442_));
 sky130_fd_sc_hd__or2_1 _10280_ (.A(_04370_),
    .B(_04372_),
    .X(_04443_));
 sky130_fd_sc_hd__nand2_1 _10281_ (.A(_04442_),
    .B(_04443_),
    .Y(_04444_));
 sky130_fd_sc_hd__xnor2_1 _10282_ (.A(_04442_),
    .B(_04443_),
    .Y(_04445_));
 sky130_fd_sc_hd__o21ai_1 _10283_ (.A1(_04336_),
    .A2(_04337_),
    .B1(_04335_),
    .Y(_04446_));
 sky130_fd_sc_hd__nand2b_1 _10284_ (.A_N(_04445_),
    .B(_04446_),
    .Y(_04447_));
 sky130_fd_sc_hd__xnor2_1 _10285_ (.A(_04445_),
    .B(_04446_),
    .Y(_04448_));
 sky130_fd_sc_hd__o21ai_1 _10286_ (.A1(_04374_),
    .A2(_04377_),
    .B1(_04448_),
    .Y(_04449_));
 sky130_fd_sc_hd__or3_1 _10287_ (.A(_04374_),
    .B(_04377_),
    .C(_04448_),
    .X(_04450_));
 sky130_fd_sc_hd__and2_1 _10288_ (.A(_04449_),
    .B(_04450_),
    .X(_04452_));
 sky130_fd_sc_hd__or3_1 _10289_ (.A(_04308_),
    .B(_04379_),
    .C(_04380_),
    .X(_04453_));
 sky130_fd_sc_hd__nor2_1 _10290_ (.A(_04306_),
    .B(_04380_),
    .Y(_04454_));
 sky130_fd_sc_hd__o22ai_1 _10291_ (.A1(_04309_),
    .A2(_04453_),
    .B1(_04454_),
    .B2(_04379_),
    .Y(_04455_));
 sky130_fd_sc_hd__nor2_1 _10292_ (.A(_04311_),
    .B(_04453_),
    .Y(_04456_));
 sky130_fd_sc_hd__a21oi_1 _10293_ (.A1(_04138_),
    .A2(_04456_),
    .B1(_04455_),
    .Y(_04457_));
 sky130_fd_sc_hd__nand2b_1 _10294_ (.A_N(_04457_),
    .B(_04452_),
    .Y(_04458_));
 sky130_fd_sc_hd__xnor2_1 _10295_ (.A(_04452_),
    .B(_04457_),
    .Y(net112));
 sky130_fd_sc_hd__a22o_1 _10296_ (.A1(net314),
    .A2(net507),
    .B1(net501),
    .B2(net321),
    .X(_04459_));
 sky130_fd_sc_hd__nand2_1 _10297_ (.A(net314),
    .B(net501),
    .Y(_04460_));
 sky130_fd_sc_hd__and4_1 _10298_ (.A(net321),
    .B(net314),
    .C(net507),
    .D(net501),
    .X(_04462_));
 sky130_fd_sc_hd__inv_2 _10299_ (.A(_04462_),
    .Y(_04463_));
 sky130_fd_sc_hd__a31o_1 _10300_ (.A1(net314),
    .A2(net527),
    .A3(_04384_),
    .B1(_04383_),
    .X(_04464_));
 sky130_fd_sc_hd__nand4_1 _10301_ (.A(net306),
    .B(net292),
    .C(net530),
    .D(net521),
    .Y(_04465_));
 sky130_fd_sc_hd__a22o_1 _10302_ (.A1(net292),
    .A2(net530),
    .B1(net521),
    .B2(net306),
    .X(_04466_));
 sky130_fd_sc_hd__nand2_1 _10303_ (.A(_04465_),
    .B(_04466_),
    .Y(_04467_));
 sky130_fd_sc_hd__nand2_1 _10304_ (.A(net284),
    .B(net537),
    .Y(_04468_));
 sky130_fd_sc_hd__xor2_1 _10305_ (.A(_04467_),
    .B(_04468_),
    .X(_04469_));
 sky130_fd_sc_hd__xor2_1 _10306_ (.A(_04464_),
    .B(_04469_),
    .X(_04470_));
 sky130_fd_sc_hd__o21ba_1 _10307_ (.A1(_04394_),
    .A2(_04397_),
    .B1_N(_04393_),
    .X(_04471_));
 sky130_fd_sc_hd__nand2b_1 _10308_ (.A_N(_04471_),
    .B(_04470_),
    .Y(_04473_));
 sky130_fd_sc_hd__xor2_1 _10309_ (.A(_04470_),
    .B(_04471_),
    .X(_04474_));
 sky130_fd_sc_hd__a21oi_1 _10310_ (.A1(_04391_),
    .A2(_04400_),
    .B1(_04399_),
    .Y(_04475_));
 sky130_fd_sc_hd__or2_1 _10311_ (.A(_04474_),
    .B(_04475_),
    .X(_04476_));
 sky130_fd_sc_hd__nand2_1 _10312_ (.A(_04474_),
    .B(_04475_),
    .Y(_04477_));
 sky130_fd_sc_hd__nand2_1 _10313_ (.A(_04476_),
    .B(_04477_),
    .Y(_04478_));
 sky130_fd_sc_hd__and2_1 _10314_ (.A(_04402_),
    .B(_04405_),
    .X(_04479_));
 sky130_fd_sc_hd__nor2_1 _10315_ (.A(_04478_),
    .B(_04479_),
    .Y(_04480_));
 sky130_fd_sc_hd__xor2_1 _10316_ (.A(_04478_),
    .B(_04479_),
    .X(_04481_));
 sky130_fd_sc_hd__and4_1 _10317_ (.A(net558),
    .B(net550),
    .C(net277),
    .D(net269),
    .X(_04482_));
 sky130_fd_sc_hd__a22oi_1 _10318_ (.A1(net550),
    .A2(net278),
    .B1(net269),
    .B2(net558),
    .Y(_04484_));
 sky130_fd_sc_hd__nor2_1 _10319_ (.A(_04482_),
    .B(_04484_),
    .Y(_04485_));
 sky130_fd_sc_hd__nand2_1 _10320_ (.A(net565),
    .B(net262),
    .Y(_04486_));
 sky130_fd_sc_hd__xnor2_1 _10321_ (.A(_04485_),
    .B(_04486_),
    .Y(_04487_));
 sky130_fd_sc_hd__o21ba_1 _10322_ (.A1(_04411_),
    .A2(_04413_),
    .B1_N(_04410_),
    .X(_04488_));
 sky130_fd_sc_hd__nand2b_1 _10323_ (.A_N(_04488_),
    .B(_04487_),
    .Y(_04489_));
 sky130_fd_sc_hd__xnor2_1 _10324_ (.A(_04487_),
    .B(_04488_),
    .Y(_04490_));
 sky130_fd_sc_hd__and2_1 _10325_ (.A(net572),
    .B(net250),
    .X(_04491_));
 sky130_fd_sc_hd__or2_1 _10326_ (.A(_04490_),
    .B(_04491_),
    .X(_04492_));
 sky130_fd_sc_hd__nand2_1 _10327_ (.A(_04490_),
    .B(_04491_),
    .Y(_04493_));
 sky130_fd_sc_hd__nand2_1 _10328_ (.A(_04492_),
    .B(_04493_),
    .Y(_04495_));
 sky130_fd_sc_hd__and3_1 _10329_ (.A(_04416_),
    .B(_04421_),
    .C(_04495_),
    .X(_04496_));
 sky130_fd_sc_hd__a21oi_1 _10330_ (.A1(_04416_),
    .A2(_04421_),
    .B1(_04495_),
    .Y(_04497_));
 sky130_fd_sc_hd__nor2_1 _10331_ (.A(_04496_),
    .B(_04497_),
    .Y(_04498_));
 sky130_fd_sc_hd__nand2_1 _10332_ (.A(net583),
    .B(net245),
    .Y(_04499_));
 sky130_fd_sc_hd__xnor2_1 _10333_ (.A(_04498_),
    .B(_04499_),
    .Y(_04500_));
 sky130_fd_sc_hd__xor2_1 _10334_ (.A(_04481_),
    .B(_04500_),
    .X(_04501_));
 sky130_fd_sc_hd__a21boi_1 _10335_ (.A1(_04408_),
    .A2(_04427_),
    .B1_N(_04409_),
    .Y(_04502_));
 sky130_fd_sc_hd__nand2b_1 _10336_ (.A_N(_04502_),
    .B(_04501_),
    .Y(_04503_));
 sky130_fd_sc_hd__xnor2_1 _10337_ (.A(_04501_),
    .B(_04502_),
    .Y(_04504_));
 sky130_fd_sc_hd__and3_1 _10338_ (.A(_04459_),
    .B(_04463_),
    .C(_04504_),
    .X(_04506_));
 sky130_fd_sc_hd__a21oi_1 _10339_ (.A1(_04459_),
    .A2(_04463_),
    .B1(_04504_),
    .Y(_04507_));
 sky130_fd_sc_hd__nor2_1 _10340_ (.A(_04506_),
    .B(_04507_),
    .Y(_04508_));
 sky130_fd_sc_hd__xor2_1 _10341_ (.A(_04436_),
    .B(_04508_),
    .X(_04509_));
 sky130_fd_sc_hd__xnor2_1 _10342_ (.A(_04434_),
    .B(_04509_),
    .Y(_04510_));
 sky130_fd_sc_hd__o21ai_1 _10343_ (.A1(_04368_),
    .A2(_04437_),
    .B1(_04439_),
    .Y(_04511_));
 sky130_fd_sc_hd__and2b_1 _10344_ (.A_N(_04510_),
    .B(_04511_),
    .X(_04512_));
 sky130_fd_sc_hd__xnor2_1 _10345_ (.A(_04510_),
    .B(_04511_),
    .Y(_04513_));
 sky130_fd_sc_hd__a32o_1 _10346_ (.A1(_04420_),
    .A2(_04421_),
    .A3(_04423_),
    .B1(_04426_),
    .B2(net585),
    .X(_04514_));
 sky130_fd_sc_hd__xnor2_1 _10347_ (.A(_04513_),
    .B(_04514_),
    .Y(_04515_));
 sky130_fd_sc_hd__nand2_1 _10348_ (.A(_04444_),
    .B(_04447_),
    .Y(_04517_));
 sky130_fd_sc_hd__a21o_1 _10349_ (.A1(_04444_),
    .A2(_04447_),
    .B1(_04515_),
    .X(_04518_));
 sky130_fd_sc_hd__and3_1 _10350_ (.A(_04444_),
    .B(_04447_),
    .C(_04515_),
    .X(_04519_));
 sky130_fd_sc_hd__xnor2_1 _10351_ (.A(_04515_),
    .B(_04517_),
    .Y(_04520_));
 sky130_fd_sc_hd__nand2_1 _10352_ (.A(_04449_),
    .B(_04458_),
    .Y(_04521_));
 sky130_fd_sc_hd__xor2_1 _10353_ (.A(_04520_),
    .B(_04521_),
    .X(net113));
 sky130_fd_sc_hd__and2_1 _10354_ (.A(net291),
    .B(net507),
    .X(_04522_));
 sky130_fd_sc_hd__nand2_1 _10355_ (.A(net291),
    .B(net507),
    .Y(_04523_));
 sky130_fd_sc_hd__and3_1 _10356_ (.A(net306),
    .B(net528),
    .C(_04522_),
    .X(_04524_));
 sky130_fd_sc_hd__a22oi_1 _10357_ (.A1(net292),
    .A2(net528),
    .B1(net507),
    .B2(net306),
    .Y(_04525_));
 sky130_fd_sc_hd__o2bb2a_1 _10358_ (.A1_N(net284),
    .A2_N(net530),
    .B1(_04524_),
    .B2(_04525_),
    .X(_04527_));
 sky130_fd_sc_hd__and4bb_1 _10359_ (.A_N(_04524_),
    .B_N(_04525_),
    .C(net284),
    .D(net530),
    .X(_04528_));
 sky130_fd_sc_hd__nor2_1 _10360_ (.A(_04527_),
    .B(_04528_),
    .Y(_04529_));
 sky130_fd_sc_hd__xnor2_1 _10361_ (.A(_04462_),
    .B(_04529_),
    .Y(_04530_));
 sky130_fd_sc_hd__o21ai_1 _10362_ (.A1(_04467_),
    .A2(_04468_),
    .B1(_04465_),
    .Y(_04531_));
 sky130_fd_sc_hd__and2b_1 _10363_ (.A_N(_04530_),
    .B(_04531_),
    .X(_04532_));
 sky130_fd_sc_hd__xor2_1 _10364_ (.A(_04530_),
    .B(_04531_),
    .X(_04533_));
 sky130_fd_sc_hd__a21bo_1 _10365_ (.A1(_04464_),
    .A2(_04469_),
    .B1_N(_04473_),
    .X(_04534_));
 sky130_fd_sc_hd__and2b_1 _10366_ (.A_N(_04533_),
    .B(_04534_),
    .X(_04535_));
 sky130_fd_sc_hd__xor2_1 _10367_ (.A(_04533_),
    .B(_04534_),
    .X(_04536_));
 sky130_fd_sc_hd__and2_1 _10368_ (.A(_04476_),
    .B(_04536_),
    .X(_04538_));
 sky130_fd_sc_hd__nor2_1 _10369_ (.A(_04476_),
    .B(_04536_),
    .Y(_04539_));
 sky130_fd_sc_hd__nor2_1 _10370_ (.A(_04538_),
    .B(_04539_),
    .Y(_04540_));
 sky130_fd_sc_hd__and4_1 _10371_ (.A(net551),
    .B(net537),
    .C(net277),
    .D(net269),
    .X(_04541_));
 sky130_fd_sc_hd__a22oi_1 _10372_ (.A1(net537),
    .A2(net278),
    .B1(net269),
    .B2(net551),
    .Y(_04542_));
 sky130_fd_sc_hd__nor2_1 _10373_ (.A(_04541_),
    .B(_04542_),
    .Y(_04543_));
 sky130_fd_sc_hd__nand2_1 _10374_ (.A(net558),
    .B(net262),
    .Y(_04544_));
 sky130_fd_sc_hd__xnor2_1 _10375_ (.A(_04543_),
    .B(_04544_),
    .Y(_04545_));
 sky130_fd_sc_hd__o21ba_1 _10376_ (.A1(_04484_),
    .A2(_04486_),
    .B1_N(_04482_),
    .X(_04546_));
 sky130_fd_sc_hd__nand2b_1 _10377_ (.A_N(_04546_),
    .B(_04545_),
    .Y(_04547_));
 sky130_fd_sc_hd__xnor2_1 _10378_ (.A(_04545_),
    .B(_04546_),
    .Y(_04549_));
 sky130_fd_sc_hd__and2_1 _10379_ (.A(net565),
    .B(net250),
    .X(_04550_));
 sky130_fd_sc_hd__or2_1 _10380_ (.A(_04549_),
    .B(_04550_),
    .X(_04551_));
 sky130_fd_sc_hd__nand2_1 _10381_ (.A(_04549_),
    .B(_04550_),
    .Y(_04552_));
 sky130_fd_sc_hd__nand2_1 _10382_ (.A(_04551_),
    .B(_04552_),
    .Y(_04553_));
 sky130_fd_sc_hd__and3_1 _10383_ (.A(_04489_),
    .B(_04493_),
    .C(_04553_),
    .X(_04554_));
 sky130_fd_sc_hd__a21oi_1 _10384_ (.A1(_04489_),
    .A2(_04493_),
    .B1(_04553_),
    .Y(_04555_));
 sky130_fd_sc_hd__nor2_1 _10385_ (.A(_04554_),
    .B(_04555_),
    .Y(_04556_));
 sky130_fd_sc_hd__nand2_1 _10386_ (.A(net572),
    .B(net245),
    .Y(_04557_));
 sky130_fd_sc_hd__xnor2_1 _10387_ (.A(_04556_),
    .B(_04557_),
    .Y(_04558_));
 sky130_fd_sc_hd__xnor2_1 _10388_ (.A(_04540_),
    .B(_04558_),
    .Y(_04560_));
 sky130_fd_sc_hd__a21oi_2 _10389_ (.A1(_04481_),
    .A2(_04500_),
    .B1(_04480_),
    .Y(_04561_));
 sky130_fd_sc_hd__xnor2_1 _10390_ (.A(_04560_),
    .B(_04561_),
    .Y(_04562_));
 sky130_fd_sc_hd__nor2_1 _10391_ (.A(_04460_),
    .B(_04562_),
    .Y(_04563_));
 sky130_fd_sc_hd__xor2_1 _10392_ (.A(_04460_),
    .B(_04562_),
    .X(_04564_));
 sky130_fd_sc_hd__nand2_1 _10393_ (.A(_04506_),
    .B(_04564_),
    .Y(_04565_));
 sky130_fd_sc_hd__xnor2_1 _10394_ (.A(_04506_),
    .B(_04564_),
    .Y(_04566_));
 sky130_fd_sc_hd__xnor2_1 _10395_ (.A(_04503_),
    .B(_04566_),
    .Y(_04567_));
 sky130_fd_sc_hd__o21ai_1 _10396_ (.A1(_04434_),
    .A2(_04436_),
    .B1(_04508_),
    .Y(_04568_));
 sky130_fd_sc_hd__or2_1 _10397_ (.A(_04567_),
    .B(_04568_),
    .X(_04569_));
 sky130_fd_sc_hd__xnor2_1 _10398_ (.A(_04567_),
    .B(_04568_),
    .Y(_04571_));
 sky130_fd_sc_hd__o21ba_1 _10399_ (.A1(_04496_),
    .A2(_04499_),
    .B1_N(_04497_),
    .X(_04572_));
 sky130_fd_sc_hd__or2_1 _10400_ (.A(_04571_),
    .B(_04572_),
    .X(_04573_));
 sky130_fd_sc_hd__nand2_1 _10401_ (.A(_04571_),
    .B(_04572_),
    .Y(_04574_));
 sky130_fd_sc_hd__nand2_1 _10402_ (.A(_04573_),
    .B(_04574_),
    .Y(_04575_));
 sky130_fd_sc_hd__a21oi_1 _10403_ (.A1(_04513_),
    .A2(_04514_),
    .B1(_04512_),
    .Y(_04576_));
 sky130_fd_sc_hd__nor2_1 _10404_ (.A(_04575_),
    .B(_04576_),
    .Y(_04577_));
 sky130_fd_sc_hd__or2_1 _10405_ (.A(_04575_),
    .B(_04576_),
    .X(_04578_));
 sky130_fd_sc_hd__and2_1 _10406_ (.A(_04575_),
    .B(_04576_),
    .X(_04579_));
 sky130_fd_sc_hd__nor2_1 _10407_ (.A(_04577_),
    .B(_04579_),
    .Y(_04580_));
 sky130_fd_sc_hd__a21o_1 _10408_ (.A1(_04449_),
    .A2(_04518_),
    .B1(_04519_),
    .X(_04582_));
 sky130_fd_sc_hd__nand2_1 _10409_ (.A(_04452_),
    .B(_04520_),
    .Y(_04583_));
 sky130_fd_sc_hd__o21a_1 _10410_ (.A1(_04457_),
    .A2(_04583_),
    .B1(_04582_),
    .X(_04584_));
 sky130_fd_sc_hd__xnor2_1 _10411_ (.A(_04580_),
    .B(_04584_),
    .Y(net114));
 sky130_fd_sc_hd__o21ai_1 _10412_ (.A1(_04503_),
    .A2(_04566_),
    .B1(_04565_),
    .Y(_04585_));
 sky130_fd_sc_hd__a21oi_1 _10413_ (.A1(net306),
    .A2(net501),
    .B1(_04522_),
    .Y(_04586_));
 sky130_fd_sc_hd__and3_1 _10414_ (.A(net306),
    .B(net501),
    .C(_04522_),
    .X(_04587_));
 sky130_fd_sc_hd__nor2_1 _10415_ (.A(_04586_),
    .B(_04587_),
    .Y(_04588_));
 sky130_fd_sc_hd__nand2_1 _10416_ (.A(net285),
    .B(net528),
    .Y(_04589_));
 sky130_fd_sc_hd__xnor2_1 _10417_ (.A(_04588_),
    .B(_04589_),
    .Y(_04590_));
 sky130_fd_sc_hd__o21a_1 _10418_ (.A1(_04524_),
    .A2(_04528_),
    .B1(_04590_),
    .X(_04592_));
 sky130_fd_sc_hd__nor3_1 _10419_ (.A(_04524_),
    .B(_04528_),
    .C(_04590_),
    .Y(_04593_));
 sky130_fd_sc_hd__or2_1 _10420_ (.A(_04592_),
    .B(_04593_),
    .X(_04594_));
 sky130_fd_sc_hd__a21oi_1 _10421_ (.A1(_04462_),
    .A2(_04529_),
    .B1(_04532_),
    .Y(_04595_));
 sky130_fd_sc_hd__nor2_1 _10422_ (.A(_04594_),
    .B(_04595_),
    .Y(_04596_));
 sky130_fd_sc_hd__and2_1 _10423_ (.A(_04594_),
    .B(_04595_),
    .X(_04597_));
 sky130_fd_sc_hd__nor2_1 _10424_ (.A(_04596_),
    .B(_04597_),
    .Y(_04598_));
 sky130_fd_sc_hd__xnor2_1 _10425_ (.A(_04535_),
    .B(_04598_),
    .Y(_04599_));
 sky130_fd_sc_hd__and4_1 _10426_ (.A(net536),
    .B(net279),
    .C(net529),
    .D(net271),
    .X(_04600_));
 sky130_fd_sc_hd__a22oi_1 _10427_ (.A1(net279),
    .A2(net529),
    .B1(net271),
    .B2(net536),
    .Y(_04601_));
 sky130_fd_sc_hd__nor2_1 _10428_ (.A(_04600_),
    .B(_04601_),
    .Y(_04603_));
 sky130_fd_sc_hd__nand2_1 _10429_ (.A(net551),
    .B(net261),
    .Y(_04604_));
 sky130_fd_sc_hd__xnor2_1 _10430_ (.A(_04603_),
    .B(_04604_),
    .Y(_04605_));
 sky130_fd_sc_hd__o21ba_1 _10431_ (.A1(_04542_),
    .A2(_04544_),
    .B1_N(_04541_),
    .X(_04606_));
 sky130_fd_sc_hd__nand2b_1 _10432_ (.A_N(_04606_),
    .B(_04605_),
    .Y(_04607_));
 sky130_fd_sc_hd__xnor2_1 _10433_ (.A(_04605_),
    .B(_04606_),
    .Y(_04608_));
 sky130_fd_sc_hd__and2_1 _10434_ (.A(net558),
    .B(net250),
    .X(_04609_));
 sky130_fd_sc_hd__or2_1 _10435_ (.A(_04608_),
    .B(_04609_),
    .X(_04610_));
 sky130_fd_sc_hd__nand2_1 _10436_ (.A(_04608_),
    .B(_04609_),
    .Y(_04611_));
 sky130_fd_sc_hd__nand2_1 _10437_ (.A(_04610_),
    .B(_04611_),
    .Y(_04612_));
 sky130_fd_sc_hd__and3_1 _10438_ (.A(_04547_),
    .B(_04552_),
    .C(_04612_),
    .X(_04614_));
 sky130_fd_sc_hd__a21oi_1 _10439_ (.A1(_04547_),
    .A2(_04552_),
    .B1(_04612_),
    .Y(_04615_));
 sky130_fd_sc_hd__nor2_1 _10440_ (.A(_04614_),
    .B(_04615_),
    .Y(_04616_));
 sky130_fd_sc_hd__nand2_1 _10441_ (.A(net565),
    .B(net245),
    .Y(_04617_));
 sky130_fd_sc_hd__xnor2_1 _10442_ (.A(_04616_),
    .B(_04617_),
    .Y(_04618_));
 sky130_fd_sc_hd__and2b_1 _10443_ (.A_N(_04599_),
    .B(_04618_),
    .X(_04619_));
 sky130_fd_sc_hd__xnor2_1 _10444_ (.A(_04599_),
    .B(_04618_),
    .Y(_04620_));
 sky130_fd_sc_hd__a21o_1 _10445_ (.A1(_04540_),
    .A2(_04558_),
    .B1(_04539_),
    .X(_04621_));
 sky130_fd_sc_hd__and2_1 _10446_ (.A(_04620_),
    .B(_04621_),
    .X(_04622_));
 sky130_fd_sc_hd__nor2_1 _10447_ (.A(_04620_),
    .B(_04621_),
    .Y(_04623_));
 sky130_fd_sc_hd__nor2_1 _10448_ (.A(_04622_),
    .B(_04623_),
    .Y(_04625_));
 sky130_fd_sc_hd__o21bai_2 _10449_ (.A1(_04560_),
    .A2(_04561_),
    .B1_N(_04563_),
    .Y(_04626_));
 sky130_fd_sc_hd__xor2_1 _10450_ (.A(_04625_),
    .B(_04626_),
    .X(_04627_));
 sky130_fd_sc_hd__nand2_1 _10451_ (.A(_04585_),
    .B(_04627_),
    .Y(_04628_));
 sky130_fd_sc_hd__xnor2_1 _10452_ (.A(_04585_),
    .B(_04627_),
    .Y(_04629_));
 sky130_fd_sc_hd__o21ba_1 _10453_ (.A1(_04554_),
    .A2(_04557_),
    .B1_N(_04555_),
    .X(_04630_));
 sky130_fd_sc_hd__xnor2_1 _10454_ (.A(_04629_),
    .B(_04630_),
    .Y(_04631_));
 sky130_fd_sc_hd__and3_1 _10455_ (.A(_04569_),
    .B(_04573_),
    .C(_04631_),
    .X(_04632_));
 sky130_fd_sc_hd__a21o_1 _10456_ (.A1(_04569_),
    .A2(_04573_),
    .B1(_04631_),
    .X(_04633_));
 sky130_fd_sc_hd__and2b_1 _10457_ (.A_N(_04632_),
    .B(_04633_),
    .X(_04634_));
 sky130_fd_sc_hd__o21ai_1 _10458_ (.A1(_04579_),
    .A2(_04584_),
    .B1(_04578_),
    .Y(_04636_));
 sky130_fd_sc_hd__xor2_1 _10459_ (.A(_04634_),
    .B(_04636_),
    .X(net115));
 sky130_fd_sc_hd__a31o_1 _10460_ (.A1(net565),
    .A2(net245),
    .A3(_04616_),
    .B1(_04615_),
    .X(_04637_));
 sky130_fd_sc_hd__and4_1 _10461_ (.A(net279),
    .B(net529),
    .C(net271),
    .D(net521),
    .X(_04638_));
 sky130_fd_sc_hd__a22oi_1 _10462_ (.A1(net529),
    .A2(net271),
    .B1(net521),
    .B2(net279),
    .Y(_04639_));
 sky130_fd_sc_hd__nor2_1 _10463_ (.A(_04638_),
    .B(_04639_),
    .Y(_04640_));
 sky130_fd_sc_hd__nand2_1 _10464_ (.A(net536),
    .B(net261),
    .Y(_04641_));
 sky130_fd_sc_hd__xnor2_1 _10465_ (.A(_04640_),
    .B(_04641_),
    .Y(_04642_));
 sky130_fd_sc_hd__o21ba_1 _10466_ (.A1(_04601_),
    .A2(_04604_),
    .B1_N(_04600_),
    .X(_04643_));
 sky130_fd_sc_hd__nand2b_1 _10467_ (.A_N(_04643_),
    .B(_04642_),
    .Y(_04644_));
 sky130_fd_sc_hd__xnor2_1 _10468_ (.A(_04642_),
    .B(_04643_),
    .Y(_04646_));
 sky130_fd_sc_hd__and2_1 _10469_ (.A(net551),
    .B(net251),
    .X(_04647_));
 sky130_fd_sc_hd__or2_1 _10470_ (.A(_04646_),
    .B(_04647_),
    .X(_04648_));
 sky130_fd_sc_hd__nand2_1 _10471_ (.A(_04646_),
    .B(_04647_),
    .Y(_04649_));
 sky130_fd_sc_hd__nand2_1 _10472_ (.A(_04648_),
    .B(_04649_),
    .Y(_04650_));
 sky130_fd_sc_hd__and3_1 _10473_ (.A(_04607_),
    .B(_04611_),
    .C(_04650_),
    .X(_04651_));
 sky130_fd_sc_hd__a21oi_1 _10474_ (.A1(_04607_),
    .A2(_04611_),
    .B1(_04650_),
    .Y(_04652_));
 sky130_fd_sc_hd__nor2_1 _10475_ (.A(_04651_),
    .B(_04652_),
    .Y(_04653_));
 sky130_fd_sc_hd__nand2_1 _10476_ (.A(net558),
    .B(net244),
    .Y(_04654_));
 sky130_fd_sc_hd__xnor2_1 _10477_ (.A(_04653_),
    .B(_04654_),
    .Y(_04655_));
 sky130_fd_sc_hd__a31o_1 _10478_ (.A1(net285),
    .A2(net528),
    .A3(_04588_),
    .B1(_04587_),
    .X(_04657_));
 sky130_fd_sc_hd__a22oi_1 _10479_ (.A1(net284),
    .A2(net507),
    .B1(net501),
    .B2(net291),
    .Y(_04658_));
 sky130_fd_sc_hd__and4_1 _10480_ (.A(net291),
    .B(net284),
    .C(net507),
    .D(net25),
    .X(_04659_));
 sky130_fd_sc_hd__nor2_1 _10481_ (.A(_04658_),
    .B(_04659_),
    .Y(_04660_));
 sky130_fd_sc_hd__nand2_1 _10482_ (.A(_04657_),
    .B(_04660_),
    .Y(_04661_));
 sky130_fd_sc_hd__xor2_2 _10483_ (.A(_04657_),
    .B(_04660_),
    .X(_04662_));
 sky130_fd_sc_hd__nor2_1 _10484_ (.A(_04592_),
    .B(_04596_),
    .Y(_04663_));
 sky130_fd_sc_hd__xnor2_1 _10485_ (.A(_04662_),
    .B(_04663_),
    .Y(_04664_));
 sky130_fd_sc_hd__xor2_1 _10486_ (.A(_04655_),
    .B(_04664_),
    .X(_04665_));
 sky130_fd_sc_hd__a21o_1 _10487_ (.A1(_04535_),
    .A2(_04598_),
    .B1(_04619_),
    .X(_04666_));
 sky130_fd_sc_hd__and2_1 _10488_ (.A(_04665_),
    .B(_04666_),
    .X(_04668_));
 sky130_fd_sc_hd__nor2_1 _10489_ (.A(_04665_),
    .B(_04666_),
    .Y(_04669_));
 sky130_fd_sc_hd__nor2_1 _10490_ (.A(_04668_),
    .B(_04669_),
    .Y(_04670_));
 sky130_fd_sc_hd__a21o_1 _10491_ (.A1(_04625_),
    .A2(_04626_),
    .B1(_04622_),
    .X(_04671_));
 sky130_fd_sc_hd__and2_1 _10492_ (.A(_04622_),
    .B(_04670_),
    .X(_04672_));
 sky130_fd_sc_hd__and3_1 _10493_ (.A(_04625_),
    .B(_04626_),
    .C(_04670_),
    .X(_04673_));
 sky130_fd_sc_hd__xnor2_1 _10494_ (.A(_04670_),
    .B(_04671_),
    .Y(_04674_));
 sky130_fd_sc_hd__and2b_1 _10495_ (.A_N(_04674_),
    .B(_04637_),
    .X(_04675_));
 sky130_fd_sc_hd__xor2_1 _10496_ (.A(_04637_),
    .B(_04674_),
    .X(_04676_));
 sky130_fd_sc_hd__o21a_1 _10497_ (.A1(_04629_),
    .A2(_04630_),
    .B1(_04628_),
    .X(_04677_));
 sky130_fd_sc_hd__nor2_1 _10498_ (.A(_04676_),
    .B(_04677_),
    .Y(_04679_));
 sky130_fd_sc_hd__and2_1 _10499_ (.A(_04676_),
    .B(_04677_),
    .X(_04680_));
 sky130_fd_sc_hd__nor2_1 _10500_ (.A(_04679_),
    .B(_04680_),
    .Y(_04681_));
 sky130_fd_sc_hd__nand2_1 _10501_ (.A(_04580_),
    .B(_04634_),
    .Y(_04682_));
 sky130_fd_sc_hd__nor2_1 _10502_ (.A(_04583_),
    .B(_04682_),
    .Y(_04683_));
 sky130_fd_sc_hd__a21oi_1 _10503_ (.A1(_04578_),
    .A2(_04633_),
    .B1(_04632_),
    .Y(_04684_));
 sky130_fd_sc_hd__a2bb2o_1 _10504_ (.A1_N(_04582_),
    .A2_N(_04682_),
    .B1(_04683_),
    .B2(_04455_),
    .X(_04685_));
 sky130_fd_sc_hd__a311o_1 _10505_ (.A1(_04138_),
    .A2(_04456_),
    .A3(_04683_),
    .B1(_04684_),
    .C1(_04685_),
    .X(_04686_));
 sky130_fd_sc_hd__xor2_1 _10506_ (.A(_04681_),
    .B(_04686_),
    .X(net116));
 sky130_fd_sc_hd__a31o_1 _10507_ (.A1(net558),
    .A2(net245),
    .A3(_04653_),
    .B1(_04652_),
    .X(_04687_));
 sky130_fd_sc_hd__nand2_1 _10508_ (.A(net267),
    .B(net506),
    .Y(_04688_));
 sky130_fd_sc_hd__and4_1 _10509_ (.A(net279),
    .B(net271),
    .C(net521),
    .D(net506),
    .X(_04689_));
 sky130_fd_sc_hd__a22oi_1 _10510_ (.A1(net271),
    .A2(net521),
    .B1(net506),
    .B2(net279),
    .Y(_04690_));
 sky130_fd_sc_hd__nor2_1 _10511_ (.A(_04689_),
    .B(_04690_),
    .Y(_04691_));
 sky130_fd_sc_hd__nand2_1 _10512_ (.A(net529),
    .B(net261),
    .Y(_04692_));
 sky130_fd_sc_hd__xnor2_1 _10513_ (.A(_04691_),
    .B(_04692_),
    .Y(_04693_));
 sky130_fd_sc_hd__o21ba_1 _10514_ (.A1(_04639_),
    .A2(_04641_),
    .B1_N(_04638_),
    .X(_04694_));
 sky130_fd_sc_hd__nand2b_1 _10515_ (.A_N(_04694_),
    .B(_04693_),
    .Y(_04695_));
 sky130_fd_sc_hd__xnor2_1 _10516_ (.A(_04693_),
    .B(_04694_),
    .Y(_04696_));
 sky130_fd_sc_hd__and2_1 _10517_ (.A(net536),
    .B(net251),
    .X(_04697_));
 sky130_fd_sc_hd__or2_1 _10518_ (.A(_04696_),
    .B(_04697_),
    .X(_04699_));
 sky130_fd_sc_hd__nand2_1 _10519_ (.A(_04696_),
    .B(_04697_),
    .Y(_04700_));
 sky130_fd_sc_hd__nand2_1 _10520_ (.A(_04699_),
    .B(_04700_),
    .Y(_04701_));
 sky130_fd_sc_hd__and3_1 _10521_ (.A(_04644_),
    .B(_04649_),
    .C(_04701_),
    .X(_04702_));
 sky130_fd_sc_hd__a21oi_1 _10522_ (.A1(_04644_),
    .A2(_04649_),
    .B1(_04701_),
    .Y(_04703_));
 sky130_fd_sc_hd__nor2_1 _10523_ (.A(_04702_),
    .B(_04703_),
    .Y(_04704_));
 sky130_fd_sc_hd__nand2_1 _10524_ (.A(net551),
    .B(net244),
    .Y(_04705_));
 sky130_fd_sc_hd__xnor2_1 _10525_ (.A(_04704_),
    .B(_04705_),
    .Y(_04706_));
 sky130_fd_sc_hd__nand2_1 _10526_ (.A(net285),
    .B(net25),
    .Y(_04707_));
 sky130_fd_sc_hd__nor2_1 _10527_ (.A(_04522_),
    .B(_04707_),
    .Y(_04708_));
 sky130_fd_sc_hd__a21bo_1 _10528_ (.A1(_04592_),
    .A2(_04662_),
    .B1_N(_04661_),
    .X(_04710_));
 sky130_fd_sc_hd__xor2_1 _10529_ (.A(_04708_),
    .B(_04710_),
    .X(_04711_));
 sky130_fd_sc_hd__xor2_1 _10530_ (.A(_04706_),
    .B(_04711_),
    .X(_04712_));
 sky130_fd_sc_hd__a22o_1 _10531_ (.A1(_04596_),
    .A2(_04662_),
    .B1(_04664_),
    .B2(_04655_),
    .X(_04713_));
 sky130_fd_sc_hd__and2_1 _10532_ (.A(_04712_),
    .B(_04713_),
    .X(_04714_));
 sky130_fd_sc_hd__nor2_1 _10533_ (.A(_04712_),
    .B(_04713_),
    .Y(_04715_));
 sky130_fd_sc_hd__nor2_1 _10534_ (.A(_04714_),
    .B(_04715_),
    .Y(_04716_));
 sky130_fd_sc_hd__nand2_1 _10535_ (.A(_04668_),
    .B(_04716_),
    .Y(_04717_));
 sky130_fd_sc_hd__nand2_1 _10536_ (.A(_04672_),
    .B(_04716_),
    .Y(_04718_));
 sky130_fd_sc_hd__or3_1 _10537_ (.A(_04668_),
    .B(_04672_),
    .C(_04716_),
    .X(_04719_));
 sky130_fd_sc_hd__and3_1 _10538_ (.A(_04717_),
    .B(_04718_),
    .C(_04719_),
    .X(_04721_));
 sky130_fd_sc_hd__xor2_1 _10539_ (.A(_04687_),
    .B(_04721_),
    .X(_04722_));
 sky130_fd_sc_hd__or3_1 _10540_ (.A(_04673_),
    .B(_04675_),
    .C(_04722_),
    .X(_04723_));
 sky130_fd_sc_hd__o21ai_1 _10541_ (.A1(_04673_),
    .A2(_04675_),
    .B1(_04722_),
    .Y(_04724_));
 sky130_fd_sc_hd__and2_1 _10542_ (.A(_04723_),
    .B(_04724_),
    .X(_04725_));
 sky130_fd_sc_hd__a21oi_1 _10543_ (.A1(_04681_),
    .A2(_04686_),
    .B1(_04679_),
    .Y(_04726_));
 sky130_fd_sc_hd__xnor2_1 _10544_ (.A(_04725_),
    .B(_04726_),
    .Y(net117));
 sky130_fd_sc_hd__and4_1 _10545_ (.A(net276),
    .B(net267),
    .C(net506),
    .D(net500),
    .X(_04727_));
 sky130_fd_sc_hd__nand4_1 _10546_ (.A(net276),
    .B(net267),
    .C(net506),
    .D(net500),
    .Y(_04728_));
 sky130_fd_sc_hd__a22o_1 _10547_ (.A1(net267),
    .A2(net506),
    .B1(net500),
    .B2(net276),
    .X(_04729_));
 sky130_fd_sc_hd__and2_1 _10548_ (.A(net521),
    .B(net261),
    .X(_04731_));
 sky130_fd_sc_hd__a21oi_1 _10549_ (.A1(_04728_),
    .A2(_04729_),
    .B1(_04731_),
    .Y(_04732_));
 sky130_fd_sc_hd__and3_1 _10550_ (.A(_04728_),
    .B(_04729_),
    .C(_04731_),
    .X(_04733_));
 sky130_fd_sc_hd__nor2_1 _10551_ (.A(_04732_),
    .B(_04733_),
    .Y(_04734_));
 sky130_fd_sc_hd__o21ba_1 _10552_ (.A1(_04690_),
    .A2(_04692_),
    .B1_N(_04689_),
    .X(_04735_));
 sky130_fd_sc_hd__and2b_1 _10553_ (.A_N(_04735_),
    .B(_04734_),
    .X(_04736_));
 sky130_fd_sc_hd__xnor2_1 _10554_ (.A(_04734_),
    .B(_04735_),
    .Y(_04737_));
 sky130_fd_sc_hd__nand2_1 _10555_ (.A(net529),
    .B(net251),
    .Y(_04738_));
 sky130_fd_sc_hd__xor2_1 _10556_ (.A(_04737_),
    .B(_04738_),
    .X(_04739_));
 sky130_fd_sc_hd__and3_1 _10557_ (.A(_04695_),
    .B(_04700_),
    .C(_04739_),
    .X(_04740_));
 sky130_fd_sc_hd__a21oi_1 _10558_ (.A1(_04695_),
    .A2(_04700_),
    .B1(_04739_),
    .Y(_04742_));
 sky130_fd_sc_hd__nor2_1 _10559_ (.A(_04740_),
    .B(_04742_),
    .Y(_04743_));
 sky130_fd_sc_hd__nand2_1 _10560_ (.A(net536),
    .B(net244),
    .Y(_04744_));
 sky130_fd_sc_hd__xnor2_1 _10561_ (.A(_04743_),
    .B(_04744_),
    .Y(_04745_));
 sky130_fd_sc_hd__a21oi_1 _10562_ (.A1(_04523_),
    .A2(_04661_),
    .B1(_04707_),
    .Y(_04746_));
 sky130_fd_sc_hd__and2_1 _10563_ (.A(_04745_),
    .B(_04746_),
    .X(_04747_));
 sky130_fd_sc_hd__nor2_1 _10564_ (.A(_04745_),
    .B(_04746_),
    .Y(_04748_));
 sky130_fd_sc_hd__nor2_1 _10565_ (.A(_04747_),
    .B(_04748_),
    .Y(_04749_));
 sky130_fd_sc_hd__a32o_1 _10566_ (.A1(_04592_),
    .A2(_04662_),
    .A3(_04708_),
    .B1(_04711_),
    .B2(_04706_),
    .X(_04750_));
 sky130_fd_sc_hd__xnor2_1 _10567_ (.A(_04749_),
    .B(_04750_),
    .Y(_04751_));
 sky130_fd_sc_hd__inv_2 _10568_ (.A(_04751_),
    .Y(_04753_));
 sky130_fd_sc_hd__xnor2_1 _10569_ (.A(_04714_),
    .B(_04753_),
    .Y(_04754_));
 sky130_fd_sc_hd__or2_1 _10570_ (.A(_04717_),
    .B(_04754_),
    .X(_04755_));
 sky130_fd_sc_hd__nand2_1 _10571_ (.A(_04717_),
    .B(_04754_),
    .Y(_04756_));
 sky130_fd_sc_hd__nand2_1 _10572_ (.A(_04755_),
    .B(_04756_),
    .Y(_04757_));
 sky130_fd_sc_hd__a31o_1 _10573_ (.A1(net551),
    .A2(net244),
    .A3(_04704_),
    .B1(_04703_),
    .X(_04758_));
 sky130_fd_sc_hd__nand2b_1 _10574_ (.A_N(_04757_),
    .B(_04758_),
    .Y(_04759_));
 sky130_fd_sc_hd__xnor2_1 _10575_ (.A(_04757_),
    .B(_04758_),
    .Y(_04760_));
 sky130_fd_sc_hd__a22o_1 _10576_ (.A1(_04672_),
    .A2(_04716_),
    .B1(_04721_),
    .B2(_04687_),
    .X(_04761_));
 sky130_fd_sc_hd__and2_1 _10577_ (.A(_04760_),
    .B(_04761_),
    .X(_04762_));
 sky130_fd_sc_hd__or2_1 _10578_ (.A(_04760_),
    .B(_04761_),
    .X(_04764_));
 sky130_fd_sc_hd__and2b_1 _10579_ (.A_N(_04762_),
    .B(_04764_),
    .X(_04765_));
 sky130_fd_sc_hd__and3_1 _10580_ (.A(_04681_),
    .B(_04686_),
    .C(_04725_),
    .X(_04766_));
 sky130_fd_sc_hd__a21bo_1 _10581_ (.A1(_04679_),
    .A2(_04723_),
    .B1_N(_04724_),
    .X(_04767_));
 sky130_fd_sc_hd__o21a_1 _10582_ (.A1(_04766_),
    .A2(_04767_),
    .B1(_04765_),
    .X(_04768_));
 sky130_fd_sc_hd__nor3_1 _10583_ (.A(_04765_),
    .B(_04766_),
    .C(_04767_),
    .Y(_04769_));
 sky130_fd_sc_hd__nor2_1 _10584_ (.A(_04768_),
    .B(_04769_),
    .Y(net118));
 sky130_fd_sc_hd__nand2_1 _10585_ (.A(net260),
    .B(net500),
    .Y(_04770_));
 sky130_fd_sc_hd__a22o_1 _10586_ (.A1(net260),
    .A2(net506),
    .B1(net500),
    .B2(net267),
    .X(_04771_));
 sky130_fd_sc_hd__o21a_1 _10587_ (.A1(_04688_),
    .A2(_04770_),
    .B1(_04771_),
    .X(_04772_));
 sky130_fd_sc_hd__nor3_1 _10588_ (.A(_04727_),
    .B(_04733_),
    .C(_04772_),
    .Y(_04774_));
 sky130_fd_sc_hd__o21a_1 _10589_ (.A1(_04727_),
    .A2(_04733_),
    .B1(_04772_),
    .X(_04775_));
 sky130_fd_sc_hd__nor2_1 _10590_ (.A(_04774_),
    .B(_04775_),
    .Y(_04776_));
 sky130_fd_sc_hd__nand2_1 _10591_ (.A(net521),
    .B(net249),
    .Y(_04777_));
 sky130_fd_sc_hd__xor2_1 _10592_ (.A(_04776_),
    .B(_04777_),
    .X(_04778_));
 sky130_fd_sc_hd__a31oi_2 _10593_ (.A1(net529),
    .A2(net251),
    .A3(_04737_),
    .B1(_04736_),
    .Y(_04779_));
 sky130_fd_sc_hd__xnor2_1 _10594_ (.A(_04778_),
    .B(_04779_),
    .Y(_04780_));
 sky130_fd_sc_hd__nand2_1 _10595_ (.A(net529),
    .B(net243),
    .Y(_04781_));
 sky130_fd_sc_hd__nor2_1 _10596_ (.A(_04780_),
    .B(_04781_),
    .Y(_04782_));
 sky130_fd_sc_hd__and2_1 _10597_ (.A(_04780_),
    .B(_04781_),
    .X(_04783_));
 sky130_fd_sc_hd__nor2_1 _10598_ (.A(_04782_),
    .B(_04783_),
    .Y(_04785_));
 sky130_fd_sc_hd__a21oi_1 _10599_ (.A1(_04749_),
    .A2(_04750_),
    .B1(_04747_),
    .Y(_04786_));
 sky130_fd_sc_hd__nand2b_1 _10600_ (.A_N(_04786_),
    .B(_04785_),
    .Y(_04787_));
 sky130_fd_sc_hd__xnor2_1 _10601_ (.A(_04785_),
    .B(_04786_),
    .Y(_04788_));
 sky130_fd_sc_hd__and3_1 _10602_ (.A(_04714_),
    .B(_04753_),
    .C(_04788_),
    .X(_04789_));
 sky130_fd_sc_hd__a21oi_1 _10603_ (.A1(_04714_),
    .A2(_04753_),
    .B1(_04788_),
    .Y(_04790_));
 sky130_fd_sc_hd__or2_1 _10604_ (.A(_04789_),
    .B(_04790_),
    .X(_04791_));
 sky130_fd_sc_hd__o21ba_1 _10605_ (.A1(_04740_),
    .A2(_04744_),
    .B1_N(_04742_),
    .X(_04792_));
 sky130_fd_sc_hd__nor2_1 _10606_ (.A(_04791_),
    .B(_04792_),
    .Y(_04793_));
 sky130_fd_sc_hd__xnor2_1 _10607_ (.A(_04791_),
    .B(_04792_),
    .Y(_04794_));
 sky130_fd_sc_hd__nand3_1 _10608_ (.A(_04755_),
    .B(_04759_),
    .C(_04794_),
    .Y(_04796_));
 sky130_fd_sc_hd__inv_2 _10609_ (.A(_04796_),
    .Y(_04797_));
 sky130_fd_sc_hd__a21oi_1 _10610_ (.A1(_04755_),
    .A2(_04759_),
    .B1(_04794_),
    .Y(_04798_));
 sky130_fd_sc_hd__nor2_1 _10611_ (.A(_04797_),
    .B(_04798_),
    .Y(_04799_));
 sky130_fd_sc_hd__nor2_1 _10612_ (.A(_04762_),
    .B(_04768_),
    .Y(_04800_));
 sky130_fd_sc_hd__xnor2_1 _10613_ (.A(_04799_),
    .B(_04800_),
    .Y(net119));
 sky130_fd_sc_hd__o21ba_1 _10614_ (.A1(_04778_),
    .A2(_04779_),
    .B1_N(_04782_),
    .X(_04801_));
 sky130_fd_sc_hd__and3_1 _10615_ (.A(net260),
    .B(net501),
    .C(_04688_),
    .X(_04802_));
 sky130_fd_sc_hd__nand2_1 _10616_ (.A(net506),
    .B(net249),
    .Y(_04803_));
 sky130_fd_sc_hd__xor2_1 _10617_ (.A(_04802_),
    .B(_04803_),
    .X(_04804_));
 sky130_fd_sc_hd__o21ba_1 _10618_ (.A1(_04774_),
    .A2(_04777_),
    .B1_N(_04775_),
    .X(_04806_));
 sky130_fd_sc_hd__xnor2_1 _10619_ (.A(_04804_),
    .B(_04806_),
    .Y(_04807_));
 sky130_fd_sc_hd__nand2_1 _10620_ (.A(net521),
    .B(net243),
    .Y(_04808_));
 sky130_fd_sc_hd__nor2_1 _10621_ (.A(_04807_),
    .B(_04808_),
    .Y(_04809_));
 sky130_fd_sc_hd__and2_1 _10622_ (.A(_04807_),
    .B(_04808_),
    .X(_04810_));
 sky130_fd_sc_hd__nor2_1 _10623_ (.A(_04809_),
    .B(_04810_),
    .Y(_04811_));
 sky130_fd_sc_hd__xnor2_1 _10624_ (.A(_04787_),
    .B(_04811_),
    .Y(_04812_));
 sky130_fd_sc_hd__and2b_1 _10625_ (.A_N(_04801_),
    .B(_04812_),
    .X(_04813_));
 sky130_fd_sc_hd__xnor2_1 _10626_ (.A(_04801_),
    .B(_04812_),
    .Y(_04814_));
 sky130_fd_sc_hd__o21a_1 _10627_ (.A1(_04789_),
    .A2(_04793_),
    .B1(_04814_),
    .X(_04815_));
 sky130_fd_sc_hd__nor3_1 _10628_ (.A(_04789_),
    .B(_04793_),
    .C(_04814_),
    .Y(_04817_));
 sky130_fd_sc_hd__or2_1 _10629_ (.A(_04815_),
    .B(_04817_),
    .X(_04818_));
 sky130_fd_sc_hd__inv_2 _10630_ (.A(_04818_),
    .Y(_04819_));
 sky130_fd_sc_hd__a31o_1 _10631_ (.A1(_04760_),
    .A2(_04761_),
    .A3(_04796_),
    .B1(_04798_),
    .X(_04820_));
 sky130_fd_sc_hd__or3_1 _10632_ (.A(_04766_),
    .B(_04767_),
    .C(_04820_),
    .X(_04821_));
 sky130_fd_sc_hd__o21a_1 _10633_ (.A1(_04764_),
    .A2(_04798_),
    .B1(_04796_),
    .X(_04822_));
 sky130_fd_sc_hd__o311a_1 _10634_ (.A1(_04766_),
    .A2(_04767_),
    .A3(_04820_),
    .B1(_04822_),
    .C1(_04819_),
    .X(_04823_));
 sky130_fd_sc_hd__a21oi_1 _10635_ (.A1(_04821_),
    .A2(_04822_),
    .B1(_04819_),
    .Y(_04824_));
 sky130_fd_sc_hd__nor2_1 _10636_ (.A(_04823_),
    .B(_04824_),
    .Y(net121));
 sky130_fd_sc_hd__and2_1 _10637_ (.A(_04785_),
    .B(_04811_),
    .X(_04825_));
 sky130_fd_sc_hd__a21oi_1 _10638_ (.A1(_04688_),
    .A2(_04803_),
    .B1(_04770_),
    .Y(_04827_));
 sky130_fd_sc_hd__a21oi_1 _10639_ (.A1(net249),
    .A2(net500),
    .B1(_04827_),
    .Y(_04828_));
 sky130_fd_sc_hd__a41o_1 _10640_ (.A1(net260),
    .A2(net506),
    .A3(net249),
    .A4(net500),
    .B1(_04828_),
    .X(_04829_));
 sky130_fd_sc_hd__nand2_1 _10641_ (.A(net506),
    .B(net243),
    .Y(_04830_));
 sky130_fd_sc_hd__nor2_1 _10642_ (.A(_04829_),
    .B(_04830_),
    .Y(_04831_));
 sky130_fd_sc_hd__and2_1 _10643_ (.A(_04829_),
    .B(_04830_),
    .X(_04832_));
 sky130_fd_sc_hd__nor2_1 _10644_ (.A(_04831_),
    .B(_04832_),
    .Y(_04833_));
 sky130_fd_sc_hd__a21oi_1 _10645_ (.A1(_04747_),
    .A2(_04825_),
    .B1(_04833_),
    .Y(_04834_));
 sky130_fd_sc_hd__and3_1 _10646_ (.A(_04747_),
    .B(_04825_),
    .C(_04833_),
    .X(_04835_));
 sky130_fd_sc_hd__nor2_1 _10647_ (.A(_04834_),
    .B(_04835_),
    .Y(_04836_));
 sky130_fd_sc_hd__o21ba_1 _10648_ (.A1(_04804_),
    .A2(_04806_),
    .B1_N(_04809_),
    .X(_04838_));
 sky130_fd_sc_hd__and2b_1 _10649_ (.A_N(_04838_),
    .B(_04836_),
    .X(_04839_));
 sky130_fd_sc_hd__xnor2_1 _10650_ (.A(_04836_),
    .B(_04838_),
    .Y(_04840_));
 sky130_fd_sc_hd__and3_1 _10651_ (.A(_04749_),
    .B(_04750_),
    .C(_04825_),
    .X(_04841_));
 sky130_fd_sc_hd__nor3_1 _10652_ (.A(_04813_),
    .B(_04840_),
    .C(_04841_),
    .Y(_04842_));
 sky130_fd_sc_hd__o21a_1 _10653_ (.A1(_04813_),
    .A2(_04841_),
    .B1(_04840_),
    .X(_04843_));
 sky130_fd_sc_hd__nor2_1 _10654_ (.A(_04842_),
    .B(_04843_),
    .Y(_04844_));
 sky130_fd_sc_hd__nor2_1 _10655_ (.A(_04815_),
    .B(_04823_),
    .Y(_04845_));
 sky130_fd_sc_hd__xnor2_1 _10656_ (.A(_04844_),
    .B(_04845_),
    .Y(net122));
 sky130_fd_sc_hd__a31o_1 _10657_ (.A1(net249),
    .A2(net500),
    .A3(_04827_),
    .B1(_04831_),
    .X(_04846_));
 sky130_fd_sc_hd__and3_1 _10658_ (.A(net500),
    .B(net243),
    .C(_04846_),
    .X(_04848_));
 sky130_fd_sc_hd__a21oi_1 _10659_ (.A1(net500),
    .A2(net243),
    .B1(_04846_),
    .Y(_04849_));
 sky130_fd_sc_hd__or2_1 _10660_ (.A(_04848_),
    .B(_04849_),
    .X(_04850_));
 sky130_fd_sc_hd__o21ba_1 _10661_ (.A1(_04835_),
    .A2(_04839_),
    .B1_N(_04850_),
    .X(_04851_));
 sky130_fd_sc_hd__or3b_1 _10662_ (.A(_04835_),
    .B(_04839_),
    .C_N(_04850_),
    .X(_04852_));
 sky130_fd_sc_hd__nand2b_1 _10663_ (.A_N(_04851_),
    .B(_04852_),
    .Y(_04853_));
 sky130_fd_sc_hd__and2b_1 _10664_ (.A_N(_04842_),
    .B(_04815_),
    .X(_04854_));
 sky130_fd_sc_hd__a211o_1 _10665_ (.A1(_04823_),
    .A2(_04844_),
    .B1(_04854_),
    .C1(_04843_),
    .X(_04855_));
 sky130_fd_sc_hd__xnor2_1 _10666_ (.A(_04853_),
    .B(_04855_),
    .Y(net123));
 sky130_fd_sc_hd__a211o_1 _10667_ (.A1(_04852_),
    .A2(_04855_),
    .B1(_04848_),
    .C1(_04851_),
    .X(net124));
 sky130_fd_sc_hd__a21oi_1 _10668_ (.A1(_01671_),
    .A2(_02130_),
    .B1(_03255_),
    .Y(_04857_));
 sky130_fd_sc_hd__nor2_1 _10669_ (.A(_03266_),
    .B(_04857_),
    .Y(net128));
 sky130_fd_sc_hd__a22oi_1 _10670_ (.A1(net434),
    .A2(net598),
    .B1(net627),
    .B2(net341),
    .Y(_04858_));
 sky130_fd_sc_hd__nor2_1 _10671_ (.A(_00865_),
    .B(_04858_),
    .Y(net76));
 sky130_fd_sc_hd__nor2_1 _10672_ (.A(_00844_),
    .B(_00865_),
    .Y(_04859_));
 sky130_fd_sc_hd__nor2_1 _10673_ (.A(_00876_),
    .B(_04859_),
    .Y(net87));
 sky130_fd_sc_hd__nor2_1 _10674_ (.A(_00822_),
    .B(_00876_),
    .Y(_04860_));
 sky130_fd_sc_hd__nor2_1 _10675_ (.A(_00887_),
    .B(_04860_),
    .Y(net98));
 sky130_fd_sc_hd__or2_1 _10676_ (.A(_00800_),
    .B(_00887_),
    .X(_04861_));
 sky130_fd_sc_hd__and2_1 _10677_ (.A(_00898_),
    .B(_04861_),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(A[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_4 input2 (.A(A[10]),
    .X(net2));
 sky130_fd_sc_hd__buf_1 input3 (.A(A[11]),
    .X(net3));
 sky130_fd_sc_hd__buf_1 input4 (.A(A[12]),
    .X(net4));
 sky130_fd_sc_hd__buf_1 input5 (.A(A[13]),
    .X(net5));
 sky130_fd_sc_hd__buf_2 input6 (.A(A[14]),
    .X(net6));
 sky130_fd_sc_hd__buf_2 input7 (.A(A[15]),
    .X(net7));
 sky130_fd_sc_hd__buf_1 input8 (.A(A[16]),
    .X(net8));
 sky130_fd_sc_hd__buf_2 input9 (.A(A[17]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(A[18]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_2 input11 (.A(A[19]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(A[1]),
    .X(net12));
 sky130_fd_sc_hd__buf_2 input13 (.A(A[20]),
    .X(net13));
 sky130_fd_sc_hd__buf_2 input14 (.A(A[21]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(A[22]),
    .X(net15));
 sky130_fd_sc_hd__buf_2 input16 (.A(A[23]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_2 input17 (.A(A[24]),
    .X(net17));
 sky130_fd_sc_hd__buf_1 input18 (.A(A[25]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_2 input19 (.A(A[26]),
    .X(net19));
 sky130_fd_sc_hd__buf_1 input20 (.A(A[27]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_2 input21 (.A(A[28]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(A[29]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(A[2]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(A[30]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_2 input25 (.A(A[31]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_2 input26 (.A(A[3]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(A[4]),
    .X(net27));
 sky130_fd_sc_hd__buf_2 input28 (.A(A[5]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(A[6]),
    .X(net29));
 sky130_fd_sc_hd__buf_1 input30 (.A(A[7]),
    .X(net30));
 sky130_fd_sc_hd__buf_2 input31 (.A(A[8]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_4 input32 (.A(A[9]),
    .X(net32));
 sky130_fd_sc_hd__buf_1 input33 (.A(B[0]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(B[10]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(B[11]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(B[12]),
    .X(net36));
 sky130_fd_sc_hd__buf_2 input37 (.A(B[13]),
    .X(net37));
 sky130_fd_sc_hd__buf_2 input38 (.A(B[14]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_2 input39 (.A(B[15]),
    .X(net39));
 sky130_fd_sc_hd__dlymetal6s2s_1 input40 (.A(B[16]),
    .X(net40));
 sky130_fd_sc_hd__buf_1 input41 (.A(B[17]),
    .X(net41));
 sky130_fd_sc_hd__buf_2 input42 (.A(B[18]),
    .X(net42));
 sky130_fd_sc_hd__buf_2 input43 (.A(B[19]),
    .X(net43));
 sky130_fd_sc_hd__buf_2 input44 (.A(B[1]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(B[20]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_1 input46 (.A(B[21]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_2 input47 (.A(B[22]),
    .X(net47));
 sky130_fd_sc_hd__buf_2 input48 (.A(B[23]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_1 input49 (.A(B[24]),
    .X(net49));
 sky130_fd_sc_hd__buf_2 input50 (.A(B[25]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 input51 (.A(B[26]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_4 input52 (.A(B[27]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 input53 (.A(B[28]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 input54 (.A(B[29]),
    .X(net54));
 sky130_fd_sc_hd__buf_1 input55 (.A(B[2]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_1 input56 (.A(B[30]),
    .X(net56));
 sky130_fd_sc_hd__dlymetal6s2s_1 input57 (.A(B[31]),
    .X(net57));
 sky130_fd_sc_hd__buf_2 input58 (.A(B[3]),
    .X(net58));
 sky130_fd_sc_hd__buf_2 input59 (.A(B[4]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_2 input60 (.A(B[5]),
    .X(net60));
 sky130_fd_sc_hd__buf_1 input61 (.A(B[6]),
    .X(net61));
 sky130_fd_sc_hd__buf_1 input62 (.A(B[7]),
    .X(net62));
 sky130_fd_sc_hd__buf_1 input63 (.A(B[8]),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_1 input64 (.A(B[9]),
    .X(net64));
 sky130_fd_sc_hd__buf_2 output65 (.A(net65),
    .X(P[0]));
 sky130_fd_sc_hd__buf_2 output66 (.A(net66),
    .X(P[10]));
 sky130_fd_sc_hd__buf_2 output67 (.A(net67),
    .X(P[11]));
 sky130_fd_sc_hd__buf_2 output68 (.A(net68),
    .X(P[12]));
 sky130_fd_sc_hd__buf_2 output69 (.A(net69),
    .X(P[13]));
 sky130_fd_sc_hd__buf_2 output70 (.A(net70),
    .X(P[14]));
 sky130_fd_sc_hd__buf_2 output71 (.A(net71),
    .X(P[15]));
 sky130_fd_sc_hd__buf_2 output72 (.A(net72),
    .X(P[16]));
 sky130_fd_sc_hd__buf_2 output73 (.A(net73),
    .X(P[17]));
 sky130_fd_sc_hd__buf_2 output74 (.A(net74),
    .X(P[18]));
 sky130_fd_sc_hd__buf_2 output75 (.A(net75),
    .X(P[19]));
 sky130_fd_sc_hd__buf_2 output76 (.A(net76),
    .X(P[1]));
 sky130_fd_sc_hd__buf_2 output77 (.A(net77),
    .X(P[20]));
 sky130_fd_sc_hd__buf_2 output78 (.A(net78),
    .X(P[21]));
 sky130_fd_sc_hd__buf_2 output79 (.A(net79),
    .X(P[22]));
 sky130_fd_sc_hd__buf_2 output80 (.A(net80),
    .X(P[23]));
 sky130_fd_sc_hd__buf_2 output81 (.A(net81),
    .X(P[24]));
 sky130_fd_sc_hd__buf_2 output82 (.A(net82),
    .X(P[25]));
 sky130_fd_sc_hd__buf_2 output83 (.A(net83),
    .X(P[26]));
 sky130_fd_sc_hd__buf_2 output84 (.A(net84),
    .X(P[27]));
 sky130_fd_sc_hd__buf_2 output85 (.A(net85),
    .X(P[28]));
 sky130_fd_sc_hd__buf_2 output86 (.A(net86),
    .X(P[29]));
 sky130_fd_sc_hd__buf_2 output87 (.A(net87),
    .X(P[2]));
 sky130_fd_sc_hd__buf_2 output88 (.A(net88),
    .X(P[30]));
 sky130_fd_sc_hd__buf_2 output89 (.A(net89),
    .X(P[31]));
 sky130_fd_sc_hd__buf_2 output90 (.A(net90),
    .X(P[32]));
 sky130_fd_sc_hd__buf_2 output91 (.A(net91),
    .X(P[33]));
 sky130_fd_sc_hd__buf_2 output92 (.A(net92),
    .X(P[34]));
 sky130_fd_sc_hd__buf_2 output93 (.A(net93),
    .X(P[35]));
 sky130_fd_sc_hd__buf_2 output94 (.A(net94),
    .X(P[36]));
 sky130_fd_sc_hd__buf_2 output95 (.A(net95),
    .X(P[37]));
 sky130_fd_sc_hd__buf_2 output96 (.A(net96),
    .X(P[38]));
 sky130_fd_sc_hd__buf_2 output97 (.A(net97),
    .X(P[39]));
 sky130_fd_sc_hd__buf_2 output98 (.A(net98),
    .X(P[3]));
 sky130_fd_sc_hd__buf_2 output99 (.A(net99),
    .X(P[40]));
 sky130_fd_sc_hd__buf_2 output100 (.A(net100),
    .X(P[41]));
 sky130_fd_sc_hd__buf_2 output101 (.A(net101),
    .X(P[42]));
 sky130_fd_sc_hd__buf_2 output102 (.A(net102),
    .X(P[43]));
 sky130_fd_sc_hd__buf_2 output103 (.A(net103),
    .X(P[44]));
 sky130_fd_sc_hd__buf_2 output104 (.A(net104),
    .X(P[45]));
 sky130_fd_sc_hd__buf_2 output105 (.A(net105),
    .X(P[46]));
 sky130_fd_sc_hd__buf_2 output106 (.A(net106),
    .X(P[47]));
 sky130_fd_sc_hd__buf_2 output107 (.A(net107),
    .X(P[48]));
 sky130_fd_sc_hd__buf_2 output108 (.A(net108),
    .X(P[49]));
 sky130_fd_sc_hd__buf_2 output109 (.A(net109),
    .X(P[4]));
 sky130_fd_sc_hd__buf_2 output110 (.A(net110),
    .X(P[50]));
 sky130_fd_sc_hd__buf_2 output111 (.A(net111),
    .X(P[51]));
 sky130_fd_sc_hd__buf_2 output112 (.A(net112),
    .X(P[52]));
 sky130_fd_sc_hd__buf_2 output113 (.A(net113),
    .X(P[53]));
 sky130_fd_sc_hd__buf_2 output114 (.A(net114),
    .X(P[54]));
 sky130_fd_sc_hd__buf_2 output115 (.A(net115),
    .X(P[55]));
 sky130_fd_sc_hd__buf_2 output116 (.A(net116),
    .X(P[56]));
 sky130_fd_sc_hd__buf_2 output117 (.A(net117),
    .X(P[57]));
 sky130_fd_sc_hd__buf_2 output118 (.A(net118),
    .X(P[58]));
 sky130_fd_sc_hd__buf_2 output119 (.A(net119),
    .X(P[59]));
 sky130_fd_sc_hd__buf_2 output120 (.A(net120),
    .X(P[5]));
 sky130_fd_sc_hd__buf_2 output121 (.A(net121),
    .X(P[60]));
 sky130_fd_sc_hd__buf_2 output122 (.A(net122),
    .X(P[61]));
 sky130_fd_sc_hd__buf_2 output123 (.A(net123),
    .X(P[62]));
 sky130_fd_sc_hd__buf_2 output124 (.A(net124),
    .X(P[63]));
 sky130_fd_sc_hd__buf_2 output125 (.A(net125),
    .X(P[6]));
 sky130_fd_sc_hd__buf_2 output126 (.A(net126),
    .X(P[7]));
 sky130_fd_sc_hd__buf_2 output127 (.A(net127),
    .X(P[8]));
 sky130_fd_sc_hd__buf_2 output128 (.A(net128),
    .X(P[9]));
 sky130_fd_sc_hd__buf_1 max_cap129 (.A(_03120_),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_1 max_cap130 (.A(_00907_),
    .X(net130));
 sky130_fd_sc_hd__buf_1 max_cap131 (.A(_04291_),
    .X(net131));
 sky130_fd_sc_hd__buf_1 max_cap132 (.A(_01680_),
    .X(net132));
 sky130_fd_sc_hd__buf_1 max_cap133 (.A(_00902_),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_1 max_cap134 (.A(_03719_),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_1 max_cap135 (.A(_02827_),
    .X(net135));
 sky130_fd_sc_hd__buf_1 max_cap136 (.A(_04363_),
    .X(net136));
 sky130_fd_sc_hd__buf_1 max_cap137 (.A(_04204_),
    .X(net137));
 sky130_fd_sc_hd__buf_1 max_cap138 (.A(_01351_),
    .X(net138));
 sky130_fd_sc_hd__buf_1 max_cap139 (.A(_01043_),
    .X(net139));
 sky130_fd_sc_hd__buf_1 max_cap140 (.A(_01043_),
    .X(net140));
 sky130_fd_sc_hd__buf_1 max_cap141 (.A(_00749_),
    .X(net141));
 sky130_fd_sc_hd__clkbuf_1 max_cap142 (.A(_02097_),
    .X(net142));
 sky130_fd_sc_hd__clkbuf_1 max_cap143 (.A(_03061_),
    .X(net143));
 sky130_fd_sc_hd__clkbuf_1 max_cap144 (.A(_02968_),
    .X(net144));
 sky130_fd_sc_hd__clkbuf_1 wire145 (.A(_02668_),
    .X(net145));
 sky130_fd_sc_hd__clkbuf_1 max_cap146 (.A(_00893_),
    .X(net146));
 sky130_fd_sc_hd__buf_1 max_cap147 (.A(_00469_),
    .X(net147));
 sky130_fd_sc_hd__buf_1 max_cap148 (.A(_00350_),
    .X(net148));
 sky130_fd_sc_hd__buf_1 max_cap149 (.A(_00228_),
    .X(net149));
 sky130_fd_sc_hd__buf_1 max_cap150 (.A(_00125_),
    .X(net150));
 sky130_fd_sc_hd__clkbuf_1 max_cap151 (.A(_00019_),
    .X(net151));
 sky130_fd_sc_hd__clkbuf_2 max_cap152 (.A(_03323_),
    .X(net152));
 sky130_fd_sc_hd__buf_1 max_cap153 (.A(_00971_),
    .X(net153));
 sky130_fd_sc_hd__buf_1 max_cap154 (.A(_03187_),
    .X(net154));
 sky130_fd_sc_hd__buf_1 max_cap155 (.A(_02961_),
    .X(net155));
 sky130_fd_sc_hd__buf_1 max_cap156 (.A(_02775_),
    .X(net156));
 sky130_fd_sc_hd__buf_1 max_cap157 (.A(_02615_),
    .X(net157));
 sky130_fd_sc_hd__clkbuf_2 max_cap158 (.A(_01664_),
    .X(net158));
 sky130_fd_sc_hd__clkbuf_4 fanout159 (.A(net160),
    .X(net159));
 sky130_fd_sc_hd__buf_2 fanout160 (.A(net9),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_4 fanout161 (.A(net9),
    .X(net161));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout162 (.A(net9),
    .X(net162));
 sky130_fd_sc_hd__buf_2 fanout163 (.A(net166),
    .X(net163));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout164 (.A(net165),
    .X(net164));
 sky130_fd_sc_hd__buf_2 fanout165 (.A(net166),
    .X(net165));
 sky130_fd_sc_hd__buf_2 fanout166 (.A(net9),
    .X(net166));
 sky130_fd_sc_hd__buf_2 fanout167 (.A(net168),
    .X(net167));
 sky130_fd_sc_hd__clkbuf_2 fanout168 (.A(net174),
    .X(net168));
 sky130_fd_sc_hd__buf_2 fanout169 (.A(net174),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_2 fanout170 (.A(net174),
    .X(net170));
 sky130_fd_sc_hd__buf_2 fanout171 (.A(net173),
    .X(net171));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout172 (.A(net173),
    .X(net172));
 sky130_fd_sc_hd__buf_2 fanout173 (.A(net174),
    .X(net173));
 sky130_fd_sc_hd__buf_4 fanout174 (.A(net8),
    .X(net174));
 sky130_fd_sc_hd__buf_2 fanout175 (.A(net176),
    .X(net175));
 sky130_fd_sc_hd__clkbuf_2 fanout176 (.A(net7),
    .X(net176));
 sky130_fd_sc_hd__buf_2 fanout177 (.A(net7),
    .X(net177));
 sky130_fd_sc_hd__clkbuf_2 fanout178 (.A(net7),
    .X(net178));
 sky130_fd_sc_hd__buf_2 fanout179 (.A(net180),
    .X(net179));
 sky130_fd_sc_hd__buf_2 fanout180 (.A(net181),
    .X(net180));
 sky130_fd_sc_hd__clkbuf_4 fanout181 (.A(net7),
    .X(net181));
 sky130_fd_sc_hd__buf_2 fanout182 (.A(net184),
    .X(net182));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout183 (.A(net184),
    .X(net183));
 sky130_fd_sc_hd__buf_2 fanout184 (.A(net185),
    .X(net184));
 sky130_fd_sc_hd__buf_2 fanout185 (.A(net186),
    .X(net185));
 sky130_fd_sc_hd__buf_2 fanout186 (.A(net191),
    .X(net186));
 sky130_fd_sc_hd__buf_2 fanout187 (.A(net191),
    .X(net187));
 sky130_fd_sc_hd__buf_2 fanout188 (.A(net190),
    .X(net188));
 sky130_fd_sc_hd__buf_1 fanout189 (.A(net190),
    .X(net189));
 sky130_fd_sc_hd__clkbuf_2 fanout190 (.A(net191),
    .X(net190));
 sky130_fd_sc_hd__buf_2 fanout191 (.A(net64),
    .X(net191));
 sky130_fd_sc_hd__buf_2 fanout192 (.A(net194),
    .X(net192));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout193 (.A(net194),
    .X(net193));
 sky130_fd_sc_hd__clkbuf_2 fanout194 (.A(net197),
    .X(net194));
 sky130_fd_sc_hd__buf_2 fanout195 (.A(net197),
    .X(net195));
 sky130_fd_sc_hd__buf_2 fanout196 (.A(net197),
    .X(net196));
 sky130_fd_sc_hd__buf_2 fanout197 (.A(net63),
    .X(net197));
 sky130_fd_sc_hd__clkbuf_2 fanout198 (.A(net206),
    .X(net198));
 sky130_fd_sc_hd__buf_1 fanout199 (.A(net206),
    .X(net199));
 sky130_fd_sc_hd__buf_2 fanout200 (.A(net202),
    .X(net200));
 sky130_fd_sc_hd__buf_2 fanout201 (.A(net202),
    .X(net201));
 sky130_fd_sc_hd__clkbuf_2 fanout202 (.A(net206),
    .X(net202));
 sky130_fd_sc_hd__buf_2 fanout203 (.A(net205),
    .X(net203));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout204 (.A(net205),
    .X(net204));
 sky130_fd_sc_hd__buf_2 fanout205 (.A(net206),
    .X(net205));
 sky130_fd_sc_hd__buf_2 fanout206 (.A(net62),
    .X(net206));
 sky130_fd_sc_hd__clkbuf_2 fanout207 (.A(net215),
    .X(net207));
 sky130_fd_sc_hd__buf_1 fanout208 (.A(net215),
    .X(net208));
 sky130_fd_sc_hd__buf_2 fanout209 (.A(net215),
    .X(net209));
 sky130_fd_sc_hd__clkbuf_2 fanout210 (.A(net211),
    .X(net210));
 sky130_fd_sc_hd__buf_2 fanout211 (.A(net215),
    .X(net211));
 sky130_fd_sc_hd__buf_2 fanout212 (.A(net214),
    .X(net212));
 sky130_fd_sc_hd__buf_1 fanout213 (.A(net214),
    .X(net213));
 sky130_fd_sc_hd__buf_2 fanout214 (.A(net215),
    .X(net214));
 sky130_fd_sc_hd__buf_2 fanout215 (.A(net61),
    .X(net215));
 sky130_fd_sc_hd__buf_2 fanout216 (.A(net218),
    .X(net216));
 sky130_fd_sc_hd__buf_2 fanout217 (.A(net218),
    .X(net217));
 sky130_fd_sc_hd__clkbuf_4 fanout218 (.A(net60),
    .X(net218));
 sky130_fd_sc_hd__buf_2 fanout219 (.A(net60),
    .X(net219));
 sky130_fd_sc_hd__buf_2 fanout220 (.A(net223),
    .X(net220));
 sky130_fd_sc_hd__buf_2 fanout221 (.A(net223),
    .X(net221));
 sky130_fd_sc_hd__clkbuf_2 fanout222 (.A(net223),
    .X(net222));
 sky130_fd_sc_hd__buf_2 fanout223 (.A(net6),
    .X(net223));
 sky130_fd_sc_hd__buf_2 fanout224 (.A(net225),
    .X(net224));
 sky130_fd_sc_hd__buf_2 fanout225 (.A(net6),
    .X(net225));
 sky130_fd_sc_hd__buf_2 fanout226 (.A(net6),
    .X(net226));
 sky130_fd_sc_hd__clkbuf_2 fanout227 (.A(net59),
    .X(net227));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout228 (.A(net59),
    .X(net228));
 sky130_fd_sc_hd__buf_2 fanout229 (.A(net231),
    .X(net229));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout230 (.A(net231),
    .X(net230));
 sky130_fd_sc_hd__clkbuf_2 fanout231 (.A(net59),
    .X(net231));
 sky130_fd_sc_hd__clkbuf_2 fanout232 (.A(net233),
    .X(net232));
 sky130_fd_sc_hd__clkbuf_2 fanout233 (.A(net234),
    .X(net233));
 sky130_fd_sc_hd__buf_2 fanout234 (.A(net59),
    .X(net234));
 sky130_fd_sc_hd__clkbuf_2 fanout235 (.A(net58),
    .X(net235));
 sky130_fd_sc_hd__clkbuf_2 fanout236 (.A(net58),
    .X(net236));
 sky130_fd_sc_hd__clkbuf_2 fanout237 (.A(net239),
    .X(net237));
 sky130_fd_sc_hd__buf_1 fanout238 (.A(net239),
    .X(net238));
 sky130_fd_sc_hd__clkbuf_2 fanout239 (.A(net58),
    .X(net239));
 sky130_fd_sc_hd__buf_2 fanout240 (.A(net242),
    .X(net240));
 sky130_fd_sc_hd__clkbuf_2 fanout241 (.A(net242),
    .X(net241));
 sky130_fd_sc_hd__buf_2 fanout242 (.A(net58),
    .X(net242));
 sky130_fd_sc_hd__clkbuf_4 fanout243 (.A(net246),
    .X(net243));
 sky130_fd_sc_hd__clkbuf_4 fanout244 (.A(net246),
    .X(net244));
 sky130_fd_sc_hd__clkbuf_2 fanout245 (.A(net246),
    .X(net245));
 sky130_fd_sc_hd__clkbuf_4 fanout246 (.A(net57),
    .X(net246));
 sky130_fd_sc_hd__clkbuf_4 fanout247 (.A(net248),
    .X(net247));
 sky130_fd_sc_hd__buf_2 fanout248 (.A(net57),
    .X(net248));
 sky130_fd_sc_hd__clkbuf_4 fanout249 (.A(net254),
    .X(net249));
 sky130_fd_sc_hd__buf_2 fanout250 (.A(net251),
    .X(net250));
 sky130_fd_sc_hd__buf_2 fanout251 (.A(net254),
    .X(net251));
 sky130_fd_sc_hd__clkbuf_4 fanout252 (.A(net253),
    .X(net252));
 sky130_fd_sc_hd__buf_2 fanout253 (.A(net254),
    .X(net253));
 sky130_fd_sc_hd__clkbuf_4 fanout254 (.A(net56),
    .X(net254));
 sky130_fd_sc_hd__buf_2 fanout255 (.A(net258),
    .X(net255));
 sky130_fd_sc_hd__buf_2 fanout256 (.A(net257),
    .X(net256));
 sky130_fd_sc_hd__buf_2 fanout257 (.A(net258),
    .X(net257));
 sky130_fd_sc_hd__buf_2 fanout258 (.A(net55),
    .X(net258));
 sky130_fd_sc_hd__clkbuf_2 fanout259 (.A(net260),
    .X(net259));
 sky130_fd_sc_hd__buf_2 fanout260 (.A(net265),
    .X(net260));
 sky130_fd_sc_hd__buf_2 fanout261 (.A(net265),
    .X(net261));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout262 (.A(net265),
    .X(net262));
 sky130_fd_sc_hd__buf_2 fanout263 (.A(net264),
    .X(net263));
 sky130_fd_sc_hd__clkbuf_2 fanout264 (.A(net265),
    .X(net264));
 sky130_fd_sc_hd__clkbuf_4 fanout265 (.A(net54),
    .X(net265));
 sky130_fd_sc_hd__buf_2 fanout266 (.A(net268),
    .X(net266));
 sky130_fd_sc_hd__buf_1 fanout267 (.A(net268),
    .X(net267));
 sky130_fd_sc_hd__buf_2 fanout268 (.A(net274),
    .X(net268));
 sky130_fd_sc_hd__clkbuf_2 fanout269 (.A(net270),
    .X(net269));
 sky130_fd_sc_hd__buf_1 fanout270 (.A(net271),
    .X(net270));
 sky130_fd_sc_hd__buf_2 fanout271 (.A(net274),
    .X(net271));
 sky130_fd_sc_hd__buf_2 fanout272 (.A(net273),
    .X(net272));
 sky130_fd_sc_hd__clkbuf_4 fanout273 (.A(net274),
    .X(net273));
 sky130_fd_sc_hd__buf_4 fanout274 (.A(net53),
    .X(net274));
 sky130_fd_sc_hd__buf_2 fanout275 (.A(net276),
    .X(net275));
 sky130_fd_sc_hd__clkbuf_4 fanout276 (.A(net52),
    .X(net276));
 sky130_fd_sc_hd__clkbuf_2 fanout277 (.A(net278),
    .X(net277));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout278 (.A(net279),
    .X(net278));
 sky130_fd_sc_hd__clkbuf_2 fanout279 (.A(net52),
    .X(net279));
 sky130_fd_sc_hd__buf_2 fanout280 (.A(net281),
    .X(net280));
 sky130_fd_sc_hd__clkbuf_2 fanout281 (.A(net282),
    .X(net281));
 sky130_fd_sc_hd__clkbuf_4 fanout282 (.A(net52),
    .X(net282));
 sky130_fd_sc_hd__buf_4 fanout283 (.A(net286),
    .X(net283));
 sky130_fd_sc_hd__clkbuf_4 fanout284 (.A(net285),
    .X(net284));
 sky130_fd_sc_hd__clkbuf_4 fanout285 (.A(net286),
    .X(net285));
 sky130_fd_sc_hd__buf_4 fanout286 (.A(net289),
    .X(net286));
 sky130_fd_sc_hd__clkbuf_4 fanout287 (.A(net288),
    .X(net287));
 sky130_fd_sc_hd__clkbuf_4 fanout288 (.A(net289),
    .X(net288));
 sky130_fd_sc_hd__buf_2 fanout289 (.A(net51),
    .X(net289));
 sky130_fd_sc_hd__buf_4 fanout290 (.A(net293),
    .X(net290));
 sky130_fd_sc_hd__clkbuf_4 fanout291 (.A(net292),
    .X(net291));
 sky130_fd_sc_hd__clkbuf_4 fanout292 (.A(net293),
    .X(net292));
 sky130_fd_sc_hd__buf_4 fanout293 (.A(net50),
    .X(net293));
 sky130_fd_sc_hd__buf_4 fanout294 (.A(net296),
    .X(net294));
 sky130_fd_sc_hd__clkbuf_2 fanout295 (.A(net296),
    .X(net295));
 sky130_fd_sc_hd__clkbuf_4 fanout296 (.A(net50),
    .X(net296));
 sky130_fd_sc_hd__buf_2 fanout297 (.A(net299),
    .X(net297));
 sky130_fd_sc_hd__clkbuf_4 fanout298 (.A(net299),
    .X(net298));
 sky130_fd_sc_hd__clkbuf_4 fanout299 (.A(net303),
    .X(net299));
 sky130_fd_sc_hd__buf_2 fanout300 (.A(net303),
    .X(net300));
 sky130_fd_sc_hd__buf_2 fanout301 (.A(net303),
    .X(net301));
 sky130_fd_sc_hd__buf_2 fanout302 (.A(net303),
    .X(net302));
 sky130_fd_sc_hd__buf_2 fanout303 (.A(net5),
    .X(net303));
 sky130_fd_sc_hd__buf_4 fanout304 (.A(net305),
    .X(net304));
 sky130_fd_sc_hd__clkbuf_4 fanout305 (.A(net311),
    .X(net305));
 sky130_fd_sc_hd__buf_2 fanout306 (.A(net311),
    .X(net306));
 sky130_fd_sc_hd__clkbuf_4 fanout307 (.A(net311),
    .X(net307));
 sky130_fd_sc_hd__buf_4 fanout308 (.A(net311),
    .X(net308));
 sky130_fd_sc_hd__buf_2 fanout309 (.A(net311),
    .X(net309));
 sky130_fd_sc_hd__buf_2 fanout310 (.A(net311),
    .X(net310));
 sky130_fd_sc_hd__buf_4 fanout311 (.A(net49),
    .X(net311));
 sky130_fd_sc_hd__clkbuf_4 fanout312 (.A(net313),
    .X(net312));
 sky130_fd_sc_hd__clkbuf_4 fanout313 (.A(net315),
    .X(net313));
 sky130_fd_sc_hd__clkbuf_4 fanout314 (.A(net315),
    .X(net314));
 sky130_fd_sc_hd__clkbuf_2 fanout315 (.A(net48),
    .X(net315));
 sky130_fd_sc_hd__clkbuf_4 fanout316 (.A(net318),
    .X(net316));
 sky130_fd_sc_hd__clkbuf_2 fanout317 (.A(net318),
    .X(net317));
 sky130_fd_sc_hd__clkbuf_4 fanout318 (.A(net48),
    .X(net318));
 sky130_fd_sc_hd__buf_2 fanout319 (.A(net320),
    .X(net319));
 sky130_fd_sc_hd__clkbuf_4 fanout320 (.A(net322),
    .X(net320));
 sky130_fd_sc_hd__buf_2 fanout321 (.A(net322),
    .X(net321));
 sky130_fd_sc_hd__clkbuf_2 fanout322 (.A(net47),
    .X(net322));
 sky130_fd_sc_hd__clkbuf_4 fanout323 (.A(net326),
    .X(net323));
 sky130_fd_sc_hd__clkbuf_2 fanout324 (.A(net326),
    .X(net324));
 sky130_fd_sc_hd__clkbuf_4 fanout325 (.A(net326),
    .X(net325));
 sky130_fd_sc_hd__clkbuf_2 fanout326 (.A(net47),
    .X(net326));
 sky130_fd_sc_hd__buf_2 fanout327 (.A(net328),
    .X(net327));
 sky130_fd_sc_hd__clkbuf_4 fanout328 (.A(net329),
    .X(net328));
 sky130_fd_sc_hd__buf_2 fanout329 (.A(net334),
    .X(net329));
 sky130_fd_sc_hd__clkbuf_4 fanout330 (.A(net334),
    .X(net330));
 sky130_fd_sc_hd__clkbuf_2 fanout331 (.A(net334),
    .X(net331));
 sky130_fd_sc_hd__clkbuf_4 fanout332 (.A(net333),
    .X(net332));
 sky130_fd_sc_hd__clkbuf_2 fanout333 (.A(net334),
    .X(net333));
 sky130_fd_sc_hd__buf_4 fanout334 (.A(net46),
    .X(net334));
 sky130_fd_sc_hd__clkbuf_4 fanout335 (.A(net337),
    .X(net335));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout336 (.A(net337),
    .X(net336));
 sky130_fd_sc_hd__clkbuf_2 fanout337 (.A(net340),
    .X(net337));
 sky130_fd_sc_hd__clkbuf_4 fanout338 (.A(net340),
    .X(net338));
 sky130_fd_sc_hd__clkbuf_4 fanout339 (.A(net340),
    .X(net339));
 sky130_fd_sc_hd__buf_2 fanout340 (.A(net45),
    .X(net340));
 sky130_fd_sc_hd__buf_2 fanout341 (.A(net342),
    .X(net341));
 sky130_fd_sc_hd__buf_2 fanout342 (.A(net44),
    .X(net342));
 sky130_fd_sc_hd__buf_2 fanout343 (.A(net344),
    .X(net343));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout344 (.A(net348),
    .X(net344));
 sky130_fd_sc_hd__buf_2 fanout345 (.A(net346),
    .X(net345));
 sky130_fd_sc_hd__clkbuf_4 fanout346 (.A(net348),
    .X(net346));
 sky130_fd_sc_hd__buf_2 fanout347 (.A(net348),
    .X(net347));
 sky130_fd_sc_hd__buf_2 fanout348 (.A(net44),
    .X(net348));
 sky130_fd_sc_hd__buf_2 fanout349 (.A(net350),
    .X(net349));
 sky130_fd_sc_hd__clkbuf_4 fanout350 (.A(net352),
    .X(net350));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout351 (.A(net352),
    .X(net351));
 sky130_fd_sc_hd__clkbuf_4 fanout352 (.A(net43),
    .X(net352));
 sky130_fd_sc_hd__clkbuf_4 fanout353 (.A(net354),
    .X(net353));
 sky130_fd_sc_hd__buf_4 fanout354 (.A(net43),
    .X(net354));
 sky130_fd_sc_hd__buf_2 fanout355 (.A(net356),
    .X(net355));
 sky130_fd_sc_hd__clkbuf_2 fanout356 (.A(net43),
    .X(net356));
 sky130_fd_sc_hd__buf_2 fanout357 (.A(net358),
    .X(net357));
 sky130_fd_sc_hd__clkbuf_4 fanout358 (.A(net360),
    .X(net358));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout359 (.A(net360),
    .X(net359));
 sky130_fd_sc_hd__clkbuf_4 fanout360 (.A(net42),
    .X(net360));
 sky130_fd_sc_hd__clkbuf_4 fanout361 (.A(net362),
    .X(net361));
 sky130_fd_sc_hd__buf_4 fanout362 (.A(net42),
    .X(net362));
 sky130_fd_sc_hd__buf_2 fanout363 (.A(net364),
    .X(net363));
 sky130_fd_sc_hd__clkbuf_2 fanout364 (.A(net42),
    .X(net364));
 sky130_fd_sc_hd__buf_2 fanout365 (.A(net366),
    .X(net365));
 sky130_fd_sc_hd__buf_2 fanout366 (.A(net367),
    .X(net366));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout367 (.A(net372),
    .X(net367));
 sky130_fd_sc_hd__buf_2 fanout368 (.A(net369),
    .X(net368));
 sky130_fd_sc_hd__clkbuf_4 fanout369 (.A(net372),
    .X(net369));
 sky130_fd_sc_hd__clkbuf_4 fanout370 (.A(net372),
    .X(net370));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout371 (.A(net372),
    .X(net371));
 sky130_fd_sc_hd__buf_4 fanout372 (.A(net41),
    .X(net372));
 sky130_fd_sc_hd__buf_2 fanout373 (.A(net374),
    .X(net373));
 sky130_fd_sc_hd__buf_2 fanout374 (.A(net377),
    .X(net374));
 sky130_fd_sc_hd__buf_2 fanout375 (.A(net376),
    .X(net375));
 sky130_fd_sc_hd__clkbuf_4 fanout376 (.A(net377),
    .X(net376));
 sky130_fd_sc_hd__buf_2 fanout377 (.A(net40),
    .X(net377));
 sky130_fd_sc_hd__buf_2 fanout378 (.A(net380),
    .X(net378));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout379 (.A(net380),
    .X(net379));
 sky130_fd_sc_hd__clkbuf_2 fanout380 (.A(net40),
    .X(net380));
 sky130_fd_sc_hd__buf_2 fanout381 (.A(net383),
    .X(net381));
 sky130_fd_sc_hd__clkbuf_4 fanout382 (.A(net383),
    .X(net382));
 sky130_fd_sc_hd__clkbuf_4 fanout383 (.A(net388),
    .X(net383));
 sky130_fd_sc_hd__buf_2 fanout384 (.A(net388),
    .X(net384));
 sky130_fd_sc_hd__buf_1 fanout385 (.A(net388),
    .X(net385));
 sky130_fd_sc_hd__buf_2 fanout386 (.A(net388),
    .X(net386));
 sky130_fd_sc_hd__clkbuf_2 fanout387 (.A(net388),
    .X(net387));
 sky130_fd_sc_hd__buf_2 fanout388 (.A(net4),
    .X(net388));
 sky130_fd_sc_hd__buf_2 fanout389 (.A(net390),
    .X(net389));
 sky130_fd_sc_hd__buf_2 fanout390 (.A(net393),
    .X(net390));
 sky130_fd_sc_hd__buf_2 fanout391 (.A(net392),
    .X(net391));
 sky130_fd_sc_hd__clkbuf_4 fanout392 (.A(net393),
    .X(net392));
 sky130_fd_sc_hd__buf_2 fanout393 (.A(net39),
    .X(net393));
 sky130_fd_sc_hd__clkbuf_4 fanout394 (.A(net396),
    .X(net394));
 sky130_fd_sc_hd__clkbuf_2 fanout395 (.A(net396),
    .X(net395));
 sky130_fd_sc_hd__clkbuf_2 fanout396 (.A(net39),
    .X(net396));
 sky130_fd_sc_hd__clkbuf_4 fanout397 (.A(net398),
    .X(net397));
 sky130_fd_sc_hd__buf_2 fanout398 (.A(net38),
    .X(net398));
 sky130_fd_sc_hd__buf_2 fanout399 (.A(net401),
    .X(net399));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout400 (.A(net401),
    .X(net400));
 sky130_fd_sc_hd__clkbuf_2 fanout401 (.A(net38),
    .X(net401));
 sky130_fd_sc_hd__clkbuf_4 fanout402 (.A(net403),
    .X(net402));
 sky130_fd_sc_hd__buf_2 fanout403 (.A(net38),
    .X(net403));
 sky130_fd_sc_hd__clkbuf_2 fanout404 (.A(net405),
    .X(net404));
 sky130_fd_sc_hd__clkbuf_2 fanout405 (.A(net37),
    .X(net405));
 sky130_fd_sc_hd__buf_2 fanout406 (.A(net408),
    .X(net406));
 sky130_fd_sc_hd__buf_1 fanout407 (.A(net408),
    .X(net407));
 sky130_fd_sc_hd__buf_2 fanout408 (.A(net37),
    .X(net408));
 sky130_fd_sc_hd__buf_2 fanout409 (.A(net411),
    .X(net409));
 sky130_fd_sc_hd__clkbuf_2 fanout410 (.A(net411),
    .X(net410));
 sky130_fd_sc_hd__buf_2 fanout411 (.A(net37),
    .X(net411));
 sky130_fd_sc_hd__clkbuf_2 fanout412 (.A(net413),
    .X(net412));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout413 (.A(net420),
    .X(net413));
 sky130_fd_sc_hd__buf_2 fanout414 (.A(net416),
    .X(net414));
 sky130_fd_sc_hd__buf_1 fanout415 (.A(net416),
    .X(net415));
 sky130_fd_sc_hd__buf_2 fanout416 (.A(net420),
    .X(net416));
 sky130_fd_sc_hd__buf_2 fanout417 (.A(net420),
    .X(net417));
 sky130_fd_sc_hd__clkbuf_2 fanout418 (.A(net420),
    .X(net418));
 sky130_fd_sc_hd__buf_2 fanout419 (.A(net420),
    .X(net419));
 sky130_fd_sc_hd__clkbuf_4 fanout420 (.A(net36),
    .X(net420));
 sky130_fd_sc_hd__buf_2 fanout421 (.A(net422),
    .X(net421));
 sky130_fd_sc_hd__clkbuf_4 fanout422 (.A(net425),
    .X(net422));
 sky130_fd_sc_hd__buf_2 fanout423 (.A(net425),
    .X(net423));
 sky130_fd_sc_hd__clkbuf_2 fanout424 (.A(net425),
    .X(net424));
 sky130_fd_sc_hd__clkbuf_4 fanout425 (.A(net35),
    .X(net425));
 sky130_fd_sc_hd__buf_2 fanout426 (.A(net433),
    .X(net426));
 sky130_fd_sc_hd__buf_2 fanout427 (.A(net428),
    .X(net427));
 sky130_fd_sc_hd__buf_2 fanout428 (.A(net429),
    .X(net428));
 sky130_fd_sc_hd__clkbuf_2 fanout429 (.A(net433),
    .X(net429));
 sky130_fd_sc_hd__clkbuf_2 fanout430 (.A(net433),
    .X(net430));
 sky130_fd_sc_hd__buf_2 fanout431 (.A(net432),
    .X(net431));
 sky130_fd_sc_hd__buf_2 fanout432 (.A(net433),
    .X(net432));
 sky130_fd_sc_hd__clkbuf_4 fanout433 (.A(net34),
    .X(net433));
 sky130_fd_sc_hd__buf_2 fanout434 (.A(net435),
    .X(net434));
 sky130_fd_sc_hd__buf_2 fanout435 (.A(net441),
    .X(net435));
 sky130_fd_sc_hd__buf_2 fanout436 (.A(net441),
    .X(net436));
 sky130_fd_sc_hd__buf_2 fanout437 (.A(net439),
    .X(net437));
 sky130_fd_sc_hd__clkbuf_2 fanout438 (.A(net439),
    .X(net438));
 sky130_fd_sc_hd__clkbuf_2 fanout439 (.A(net441),
    .X(net439));
 sky130_fd_sc_hd__buf_2 fanout440 (.A(net441),
    .X(net440));
 sky130_fd_sc_hd__buf_2 fanout441 (.A(net33),
    .X(net441));
 sky130_fd_sc_hd__clkbuf_4 fanout442 (.A(net443),
    .X(net442));
 sky130_fd_sc_hd__buf_2 fanout443 (.A(net444),
    .X(net443));
 sky130_fd_sc_hd__buf_2 fanout444 (.A(net32),
    .X(net444));
 sky130_fd_sc_hd__buf_2 fanout445 (.A(net446),
    .X(net445));
 sky130_fd_sc_hd__clkbuf_2 fanout446 (.A(net32),
    .X(net446));
 sky130_fd_sc_hd__buf_2 fanout447 (.A(net448),
    .X(net447));
 sky130_fd_sc_hd__buf_2 fanout448 (.A(net32),
    .X(net448));
 sky130_fd_sc_hd__clkbuf_4 fanout449 (.A(net450),
    .X(net449));
 sky130_fd_sc_hd__buf_2 fanout450 (.A(net31),
    .X(net450));
 sky130_fd_sc_hd__buf_2 fanout451 (.A(net452),
    .X(net451));
 sky130_fd_sc_hd__buf_2 fanout452 (.A(net455),
    .X(net452));
 sky130_fd_sc_hd__buf_2 fanout453 (.A(net454),
    .X(net453));
 sky130_fd_sc_hd__clkbuf_2 fanout454 (.A(net455),
    .X(net454));
 sky130_fd_sc_hd__buf_2 fanout455 (.A(net31),
    .X(net455));
 sky130_fd_sc_hd__buf_2 fanout456 (.A(net457),
    .X(net456));
 sky130_fd_sc_hd__buf_2 fanout457 (.A(net462),
    .X(net457));
 sky130_fd_sc_hd__buf_2 fanout458 (.A(net459),
    .X(net458));
 sky130_fd_sc_hd__buf_2 fanout459 (.A(net462),
    .X(net459));
 sky130_fd_sc_hd__buf_2 fanout460 (.A(net462),
    .X(net460));
 sky130_fd_sc_hd__clkbuf_2 fanout461 (.A(net462),
    .X(net461));
 sky130_fd_sc_hd__buf_4 fanout462 (.A(net30),
    .X(net462));
 sky130_fd_sc_hd__clkbuf_4 fanout463 (.A(net469),
    .X(net463));
 sky130_fd_sc_hd__buf_2 fanout464 (.A(net469),
    .X(net464));
 sky130_fd_sc_hd__buf_2 fanout465 (.A(net469),
    .X(net465));
 sky130_fd_sc_hd__buf_1 fanout466 (.A(net469),
    .X(net466));
 sky130_fd_sc_hd__buf_2 fanout467 (.A(net468),
    .X(net467));
 sky130_fd_sc_hd__clkbuf_4 fanout468 (.A(net469),
    .X(net468));
 sky130_fd_sc_hd__buf_4 fanout469 (.A(net3),
    .X(net469));
 sky130_fd_sc_hd__buf_2 fanout470 (.A(net471),
    .X(net470));
 sky130_fd_sc_hd__buf_1 fanout471 (.A(net472),
    .X(net471));
 sky130_fd_sc_hd__clkbuf_2 fanout472 (.A(net477),
    .X(net472));
 sky130_fd_sc_hd__buf_2 fanout473 (.A(net474),
    .X(net473));
 sky130_fd_sc_hd__buf_2 fanout474 (.A(net477),
    .X(net474));
 sky130_fd_sc_hd__buf_2 fanout475 (.A(net477),
    .X(net475));
 sky130_fd_sc_hd__clkbuf_2 fanout476 (.A(net477),
    .X(net476));
 sky130_fd_sc_hd__clkbuf_4 fanout477 (.A(net29),
    .X(net477));
 sky130_fd_sc_hd__buf_2 fanout478 (.A(net479),
    .X(net478));
 sky130_fd_sc_hd__clkbuf_1 fanout479 (.A(net480),
    .X(net479));
 sky130_fd_sc_hd__clkbuf_2 fanout480 (.A(net28),
    .X(net480));
 sky130_fd_sc_hd__buf_2 fanout481 (.A(net482),
    .X(net481));
 sky130_fd_sc_hd__clkbuf_2 fanout482 (.A(net28),
    .X(net482));
 sky130_fd_sc_hd__buf_2 fanout483 (.A(net28),
    .X(net483));
 sky130_fd_sc_hd__clkbuf_2 fanout484 (.A(net28),
    .X(net484));
 sky130_fd_sc_hd__buf_2 fanout485 (.A(net487),
    .X(net485));
 sky130_fd_sc_hd__buf_1 fanout486 (.A(net487),
    .X(net486));
 sky130_fd_sc_hd__buf_2 fanout487 (.A(net492),
    .X(net487));
 sky130_fd_sc_hd__buf_2 fanout488 (.A(net492),
    .X(net488));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout489 (.A(net492),
    .X(net489));
 sky130_fd_sc_hd__buf_2 fanout490 (.A(net491),
    .X(net490));
 sky130_fd_sc_hd__buf_2 fanout491 (.A(net492),
    .X(net491));
 sky130_fd_sc_hd__buf_2 fanout492 (.A(net27),
    .X(net492));
 sky130_fd_sc_hd__buf_2 fanout493 (.A(net494),
    .X(net493));
 sky130_fd_sc_hd__buf_2 fanout494 (.A(net495),
    .X(net494));
 sky130_fd_sc_hd__buf_2 fanout495 (.A(net26),
    .X(net495));
 sky130_fd_sc_hd__buf_2 fanout496 (.A(net497),
    .X(net496));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout497 (.A(net26),
    .X(net497));
 sky130_fd_sc_hd__buf_2 fanout498 (.A(net499),
    .X(net498));
 sky130_fd_sc_hd__buf_2 fanout499 (.A(net26),
    .X(net499));
 sky130_fd_sc_hd__clkbuf_2 fanout500 (.A(net501),
    .X(net500));
 sky130_fd_sc_hd__clkbuf_4 fanout501 (.A(net25),
    .X(net501));
 sky130_fd_sc_hd__buf_2 fanout502 (.A(net505),
    .X(net502));
 sky130_fd_sc_hd__buf_2 fanout503 (.A(net505),
    .X(net503));
 sky130_fd_sc_hd__buf_2 fanout504 (.A(net505),
    .X(net504));
 sky130_fd_sc_hd__clkbuf_2 fanout505 (.A(net25),
    .X(net505));
 sky130_fd_sc_hd__buf_2 fanout506 (.A(net507),
    .X(net506));
 sky130_fd_sc_hd__clkbuf_4 fanout507 (.A(net24),
    .X(net507));
 sky130_fd_sc_hd__buf_2 fanout508 (.A(net513),
    .X(net508));
 sky130_fd_sc_hd__buf_2 fanout509 (.A(net510),
    .X(net509));
 sky130_fd_sc_hd__clkbuf_2 fanout510 (.A(net513),
    .X(net510));
 sky130_fd_sc_hd__buf_2 fanout511 (.A(net513),
    .X(net511));
 sky130_fd_sc_hd__clkbuf_2 fanout512 (.A(net513),
    .X(net512));
 sky130_fd_sc_hd__clkbuf_2 fanout513 (.A(net24),
    .X(net513));
 sky130_fd_sc_hd__buf_2 fanout514 (.A(net520),
    .X(net514));
 sky130_fd_sc_hd__clkbuf_2 fanout515 (.A(net520),
    .X(net515));
 sky130_fd_sc_hd__buf_2 fanout516 (.A(net520),
    .X(net516));
 sky130_fd_sc_hd__buf_2 fanout517 (.A(net520),
    .X(net517));
 sky130_fd_sc_hd__buf_2 fanout518 (.A(net519),
    .X(net518));
 sky130_fd_sc_hd__buf_2 fanout519 (.A(net520),
    .X(net519));
 sky130_fd_sc_hd__buf_4 fanout520 (.A(net23),
    .X(net520));
 sky130_fd_sc_hd__clkbuf_4 fanout521 (.A(net528),
    .X(net521));
 sky130_fd_sc_hd__buf_2 fanout522 (.A(net525),
    .X(net522));
 sky130_fd_sc_hd__buf_2 fanout523 (.A(net525),
    .X(net523));
 sky130_fd_sc_hd__clkbuf_2 fanout524 (.A(net525),
    .X(net524));
 sky130_fd_sc_hd__clkbuf_2 fanout525 (.A(net528),
    .X(net525));
 sky130_fd_sc_hd__buf_2 fanout526 (.A(net527),
    .X(net526));
 sky130_fd_sc_hd__buf_2 fanout527 (.A(net528),
    .X(net527));
 sky130_fd_sc_hd__buf_2 fanout528 (.A(net22),
    .X(net528));
 sky130_fd_sc_hd__buf_2 fanout529 (.A(net530),
    .X(net529));
 sky130_fd_sc_hd__buf_2 fanout530 (.A(net21),
    .X(net530));
 sky130_fd_sc_hd__buf_2 fanout531 (.A(net533),
    .X(net531));
 sky130_fd_sc_hd__buf_2 fanout532 (.A(net533),
    .X(net532));
 sky130_fd_sc_hd__clkbuf_2 fanout533 (.A(net21),
    .X(net533));
 sky130_fd_sc_hd__buf_2 fanout534 (.A(net535),
    .X(net534));
 sky130_fd_sc_hd__clkbuf_2 fanout535 (.A(net21),
    .X(net535));
 sky130_fd_sc_hd__buf_2 fanout536 (.A(net537),
    .X(net536));
 sky130_fd_sc_hd__buf_2 fanout537 (.A(net20),
    .X(net537));
 sky130_fd_sc_hd__buf_2 fanout538 (.A(net539),
    .X(net538));
 sky130_fd_sc_hd__buf_2 fanout539 (.A(net542),
    .X(net539));
 sky130_fd_sc_hd__buf_2 fanout540 (.A(net541),
    .X(net540));
 sky130_fd_sc_hd__buf_2 fanout541 (.A(net542),
    .X(net541));
 sky130_fd_sc_hd__clkbuf_2 fanout542 (.A(net20),
    .X(net542));
 sky130_fd_sc_hd__clkbuf_4 fanout543 (.A(net544),
    .X(net543));
 sky130_fd_sc_hd__buf_2 fanout544 (.A(net545),
    .X(net544));
 sky130_fd_sc_hd__buf_2 fanout545 (.A(net2),
    .X(net545));
 sky130_fd_sc_hd__buf_2 fanout546 (.A(net2),
    .X(net546));
 sky130_fd_sc_hd__buf_1 fanout547 (.A(net2),
    .X(net547));
 sky130_fd_sc_hd__buf_2 fanout548 (.A(net549),
    .X(net548));
 sky130_fd_sc_hd__clkbuf_4 fanout549 (.A(net2),
    .X(net549));
 sky130_fd_sc_hd__clkbuf_4 fanout550 (.A(net19),
    .X(net550));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout551 (.A(net19),
    .X(net551));
 sky130_fd_sc_hd__buf_2 fanout552 (.A(net553),
    .X(net552));
 sky130_fd_sc_hd__buf_2 fanout553 (.A(net556),
    .X(net553));
 sky130_fd_sc_hd__buf_2 fanout554 (.A(net555),
    .X(net554));
 sky130_fd_sc_hd__clkbuf_4 fanout555 (.A(net556),
    .X(net555));
 sky130_fd_sc_hd__clkbuf_2 fanout556 (.A(net19),
    .X(net556));
 sky130_fd_sc_hd__clkbuf_4 fanout557 (.A(net563),
    .X(net557));
 sky130_fd_sc_hd__clkbuf_2 fanout558 (.A(net563),
    .X(net558));
 sky130_fd_sc_hd__buf_2 fanout559 (.A(net560),
    .X(net559));
 sky130_fd_sc_hd__buf_2 fanout560 (.A(net563),
    .X(net560));
 sky130_fd_sc_hd__clkbuf_4 fanout561 (.A(net563),
    .X(net561));
 sky130_fd_sc_hd__buf_2 fanout562 (.A(net563),
    .X(net562));
 sky130_fd_sc_hd__clkbuf_4 fanout563 (.A(net18),
    .X(net563));
 sky130_fd_sc_hd__clkbuf_4 fanout564 (.A(net17),
    .X(net564));
 sky130_fd_sc_hd__clkbuf_2 fanout565 (.A(net17),
    .X(net565));
 sky130_fd_sc_hd__buf_2 fanout566 (.A(net570),
    .X(net566));
 sky130_fd_sc_hd__buf_2 fanout567 (.A(net570),
    .X(net567));
 sky130_fd_sc_hd__buf_2 fanout568 (.A(net569),
    .X(net568));
 sky130_fd_sc_hd__clkbuf_4 fanout569 (.A(net570),
    .X(net569));
 sky130_fd_sc_hd__buf_2 fanout570 (.A(net17),
    .X(net570));
 sky130_fd_sc_hd__buf_2 fanout571 (.A(net572),
    .X(net571));
 sky130_fd_sc_hd__clkbuf_4 fanout572 (.A(net16),
    .X(net572));
 sky130_fd_sc_hd__buf_2 fanout573 (.A(net574),
    .X(net573));
 sky130_fd_sc_hd__clkbuf_4 fanout574 (.A(net16),
    .X(net574));
 sky130_fd_sc_hd__buf_2 fanout575 (.A(net576),
    .X(net575));
 sky130_fd_sc_hd__clkbuf_4 fanout576 (.A(net16),
    .X(net576));
 sky130_fd_sc_hd__buf_2 fanout577 (.A(net578),
    .X(net577));
 sky130_fd_sc_hd__clkbuf_4 fanout578 (.A(net583),
    .X(net578));
 sky130_fd_sc_hd__buf_2 fanout579 (.A(net580),
    .X(net579));
 sky130_fd_sc_hd__buf_2 fanout580 (.A(net583),
    .X(net580));
 sky130_fd_sc_hd__buf_2 fanout581 (.A(net582),
    .X(net581));
 sky130_fd_sc_hd__buf_2 fanout582 (.A(net583),
    .X(net582));
 sky130_fd_sc_hd__buf_2 fanout583 (.A(net15),
    .X(net583));
 sky130_fd_sc_hd__buf_2 fanout584 (.A(net586),
    .X(net584));
 sky130_fd_sc_hd__buf_2 fanout585 (.A(net586),
    .X(net585));
 sky130_fd_sc_hd__clkbuf_4 fanout586 (.A(net14),
    .X(net586));
 sky130_fd_sc_hd__buf_2 fanout587 (.A(net588),
    .X(net587));
 sky130_fd_sc_hd__buf_2 fanout588 (.A(net14),
    .X(net588));
 sky130_fd_sc_hd__clkbuf_4 fanout589 (.A(net14),
    .X(net589));
 sky130_fd_sc_hd__buf_1 fanout590 (.A(net14),
    .X(net590));
 sky130_fd_sc_hd__buf_2 fanout591 (.A(net593),
    .X(net591));
 sky130_fd_sc_hd__buf_2 fanout592 (.A(net593),
    .X(net592));
 sky130_fd_sc_hd__buf_2 fanout593 (.A(net13),
    .X(net593));
 sky130_fd_sc_hd__buf_2 fanout594 (.A(net595),
    .X(net594));
 sky130_fd_sc_hd__clkbuf_2 fanout595 (.A(net13),
    .X(net595));
 sky130_fd_sc_hd__buf_2 fanout596 (.A(net597),
    .X(net596));
 sky130_fd_sc_hd__buf_2 fanout597 (.A(net13),
    .X(net597));
 sky130_fd_sc_hd__buf_2 fanout598 (.A(net599),
    .X(net598));
 sky130_fd_sc_hd__buf_1 fanout599 (.A(net601),
    .X(net599));
 sky130_fd_sc_hd__buf_2 fanout600 (.A(net601),
    .X(net600));
 sky130_fd_sc_hd__buf_2 fanout601 (.A(net606),
    .X(net601));
 sky130_fd_sc_hd__buf_2 fanout602 (.A(net606),
    .X(net602));
 sky130_fd_sc_hd__buf_1 fanout603 (.A(net606),
    .X(net603));
 sky130_fd_sc_hd__buf_2 fanout604 (.A(net606),
    .X(net604));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout605 (.A(net606),
    .X(net605));
 sky130_fd_sc_hd__buf_2 fanout606 (.A(net12),
    .X(net606));
 sky130_fd_sc_hd__buf_2 fanout607 (.A(net608),
    .X(net607));
 sky130_fd_sc_hd__buf_2 fanout608 (.A(net609),
    .X(net608));
 sky130_fd_sc_hd__buf_2 fanout609 (.A(net11),
    .X(net609));
 sky130_fd_sc_hd__buf_2 fanout610 (.A(net611),
    .X(net610));
 sky130_fd_sc_hd__buf_2 fanout611 (.A(net11),
    .X(net611));
 sky130_fd_sc_hd__buf_2 fanout612 (.A(net614),
    .X(net612));
 sky130_fd_sc_hd__buf_1 fanout613 (.A(net614),
    .X(net613));
 sky130_fd_sc_hd__buf_2 fanout614 (.A(net11),
    .X(net614));
 sky130_fd_sc_hd__buf_2 fanout615 (.A(net616),
    .X(net615));
 sky130_fd_sc_hd__buf_2 fanout616 (.A(net617),
    .X(net616));
 sky130_fd_sc_hd__clkbuf_2 fanout617 (.A(net10),
    .X(net617));
 sky130_fd_sc_hd__buf_2 fanout618 (.A(net619),
    .X(net618));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout619 (.A(net623),
    .X(net619));
 sky130_fd_sc_hd__buf_2 fanout620 (.A(net622),
    .X(net620));
 sky130_fd_sc_hd__buf_1 fanout621 (.A(net622),
    .X(net621));
 sky130_fd_sc_hd__buf_2 fanout622 (.A(net623),
    .X(net622));
 sky130_fd_sc_hd__clkbuf_2 fanout623 (.A(net10),
    .X(net623));
 sky130_fd_sc_hd__buf_2 fanout624 (.A(net625),
    .X(net624));
 sky130_fd_sc_hd__buf_2 fanout625 (.A(net627),
    .X(net625));
 sky130_fd_sc_hd__buf_1 fanout626 (.A(net627),
    .X(net626));
 sky130_fd_sc_hd__clkbuf_2 fanout627 (.A(net1),
    .X(net627));
 sky130_fd_sc_hd__buf_2 fanout628 (.A(net631),
    .X(net628));
 sky130_fd_sc_hd__buf_2 fanout629 (.A(net631),
    .X(net629));
 sky130_fd_sc_hd__clkbuf_2 fanout630 (.A(net631),
    .X(net630));
 sky130_fd_sc_hd__buf_2 fanout631 (.A(net1),
    .X(net631));
endmodule
